// module TestGen (input c, output reg a, b, s);
// 	wire [2:0] w;
// 	assign w = { a, b, s};
// 	initial begin
// 		$monitor($time,,, "A=%b B=%b S=%b C=%b", a, b, s, c);
// 		    { a, b, s } = 3'b000;
// 		#02 { a, b, s } = 3'b001;
// 		#02 { a, b, s } = 3'b001;
// 		#02 { a, b, s } = 3'b010;
// 		#02 { a, b, s } = 3'b011;
// 		#02 { a, b, s } = 3'b100;
// 		#02 { a, b, s } = 3'b101;
// 		#02 { a, b, s } = 3'b110;
// 		#02 { a, b, s } = 3'b111;
// 		#02 $finish;
// 	end
// endmodule

module TestGen (input [3:0] s, input c, output reg [3:0] a, b);
	wire [7:0] w;
	assign w = { a, b };
	initial begin
		$monitor($time,,, "Augend: %b Addend: %b Sum: %b Carry: %b", a, b, s, c);
			{ a, b } = 8'b00000000;
		#02 { a, b } = 8'b00000001;
		#02 { a, b } = 8'b00000010;
		#02 { a, b } = 8'b00000011;
		#02 { a, b } = 8'b00000100;
		#02 { a, b } = 8'b00000101;
		#02 { a, b } = 8'b00000110;
		#02 { a, b } = 8'b00000111;
		#02 { a, b } = 8'b00001000;
		#02 { a, b } = 8'b00001001;
		#02 { a, b } = 8'b00001010;
		#02 { a, b } = 8'b00001011;
		#02 { a, b } = 8'b00001100;
		#02 { a, b } = 8'b00001101;
		#02 { a, b } = 8'b00001110;
		#02 { a, b } = 8'b00001111;
		#02 { a, b } = 8'b00010000;
		#02 { a, b } = 8'b00010001;
		#02 { a, b } = 8'b00010010;
		#02 { a, b } = 8'b00010011;
		#02 { a, b } = 8'b00010100;
		#02 { a, b } = 8'b00010101;
		#02 { a, b } = 8'b00010110;
		#02 { a, b } = 8'b00010111;
		#02 { a, b } = 8'b00011000;
		#02 { a, b } = 8'b00011001;
		#02 { a, b } = 8'b00011010;
		#02 { a, b } = 8'b00011011;
		#02 { a, b } = 8'b00011100;
		#02 { a, b } = 8'b00011101;
		#02 { a, b } = 8'b00011110;
		#02 { a, b } = 8'b00011111;
		#02 { a, b } = 8'b00100000;
		#02 { a, b } = 8'b00100001;
		#02 { a, b } = 8'b00100010;
		#02 { a, b } = 8'b00100011;
		#02 { a, b } = 8'b00100100;
		#02 { a, b } = 8'b00100101;
		#02 { a, b } = 8'b00100110;
		#02 { a, b } = 8'b00100111;
		#02 { a, b } = 8'b00101000;
		#02 { a, b } = 8'b00101001;
		#02 { a, b } = 8'b00101010;
		#02 { a, b } = 8'b00101011;
		#02 { a, b } = 8'b00101100;
		#02 { a, b } = 8'b00101101;
		#02 { a, b } = 8'b00101110;
		#02 { a, b } = 8'b00101111;
		#02 { a, b } = 8'b00110000;
		#02 { a, b } = 8'b00110001;
		#02 { a, b } = 8'b00110010;
		#02 { a, b } = 8'b00110011;
		#02 { a, b } = 8'b00110100;
		#02 { a, b } = 8'b00110101;
		#02 { a, b } = 8'b00110110;
		#02 { a, b } = 8'b00110111;
		#02 { a, b } = 8'b00111000;
		#02 { a, b } = 8'b00111001;
		#02 { a, b } = 8'b00111010;
		#02 { a, b } = 8'b00111011;
		#02 { a, b } = 8'b00111100;
		#02 { a, b } = 8'b00111101;
		#02 { a, b } = 8'b00111110;
		#02 { a, b } = 8'b00111111;
		#02 { a, b } = 8'b01000000;
		#02 { a, b } = 8'b01000001;
		#02 { a, b } = 8'b01000010;
		#02 { a, b } = 8'b01000011;
		#02 { a, b } = 8'b01000100;
		#02 { a, b } = 8'b01000101;
		#02 { a, b } = 8'b01000110;
		#02 { a, b } = 8'b01000111;
		#02 { a, b } = 8'b01001000;
		#02 { a, b } = 8'b01001001;
		#02 { a, b } = 8'b01001010;
		#02 { a, b } = 8'b01001011;
		#02 { a, b } = 8'b01001100;
		#02 { a, b } = 8'b01001101;
		#02 { a, b } = 8'b01001110;
		#02 { a, b } = 8'b01001111;
		#02 { a, b } = 8'b01010000;
		#02 { a, b } = 8'b01010001;
		#02 { a, b } = 8'b01010010;
		#02 { a, b } = 8'b01010011;
		#02 { a, b } = 8'b01010100;
		#02 { a, b } = 8'b01010101;
		#02 { a, b } = 8'b01010110;
		#02 { a, b } = 8'b01010111;
		#02 { a, b } = 8'b01011000;
		#02 { a, b } = 8'b01011001;
		#02 { a, b } = 8'b01011010;
		#02 { a, b } = 8'b01011011;
		#02 { a, b } = 8'b01011100;
		#02 { a, b } = 8'b01011101;
		#02 { a, b } = 8'b01011110;
		#02 { a, b } = 8'b01011111;
		#02 { a, b } = 8'b01100000;
		#02 { a, b } = 8'b01100001;
		#02 { a, b } = 8'b01100010;
		#02 { a, b } = 8'b01100011;
		#02 { a, b } = 8'b01100100;
		#02 { a, b } = 8'b01100101;
		#02 { a, b } = 8'b01100110;
		#02 { a, b } = 8'b01100111;
		#02 { a, b } = 8'b01101000;
		#02 { a, b } = 8'b01101001;
		#02 { a, b } = 8'b01101010;
		#02 { a, b } = 8'b01101011;
		#02 { a, b } = 8'b01101100;
		#02 { a, b } = 8'b01101101;
		#02 { a, b } = 8'b01101110;
		#02 { a, b } = 8'b01101111;
		#02 { a, b } = 8'b01110000;
		#02 { a, b } = 8'b01110001;
		#02 { a, b } = 8'b01110010;
		#02 { a, b } = 8'b01110011;
		#02 { a, b } = 8'b01110100;
		#02 { a, b } = 8'b01110101;
		#02 { a, b } = 8'b01110110;
		#02 { a, b } = 8'b01110111;
		#02 { a, b } = 8'b01111000;
		#02 { a, b } = 8'b01111001;
		#02 { a, b } = 8'b01111010;
		#02 { a, b } = 8'b01111011;
		#02 { a, b } = 8'b01111100;
		#02 { a, b } = 8'b01111101;
		#02 { a, b } = 8'b01111110;
		#02 { a, b } = 8'b01111111;
		#02 { a, b } = 8'b10000000;
		#02 { a, b } = 8'b10000001;
		#02 { a, b } = 8'b10000010;
		#02 { a, b } = 8'b10000011;
		#02 { a, b } = 8'b10000100;
		#02 { a, b } = 8'b10000101;
		#02 { a, b } = 8'b10000110;
		#02 { a, b } = 8'b10000111;
		#02 { a, b } = 8'b10001000;
		#02 { a, b } = 8'b10001001;
		#02 { a, b } = 8'b10001010;
		#02 { a, b } = 8'b10001011;
		#02 { a, b } = 8'b10001100;
		#02 { a, b } = 8'b10001101;
		#02 { a, b } = 8'b10001110;
		#02 { a, b } = 8'b10001111;
		#02 { a, b } = 8'b10010000;
		#02 { a, b } = 8'b10010001;
		#02 { a, b } = 8'b10010010;
		#02 { a, b } = 8'b10010011;
		#02 { a, b } = 8'b10010100;
		#02 { a, b } = 8'b10010101;
		#02 { a, b } = 8'b10010110;
		#02 { a, b } = 8'b10010111;
		#02 { a, b } = 8'b10011000;
		#02 { a, b } = 8'b10011001;
		#02 { a, b } = 8'b10011010;
		#02 { a, b } = 8'b10011011;
		#02 { a, b } = 8'b10011100;
		#02 { a, b } = 8'b10011101;
		#02 { a, b } = 8'b10011110;
		#02 { a, b } = 8'b10011111;
		#02 { a, b } = 8'b10100000;
		#02 { a, b } = 8'b10100001;
		#02 { a, b } = 8'b10100010;
		#02 { a, b } = 8'b10100011;
		#02 { a, b } = 8'b10100100;
		#02 { a, b } = 8'b10100101;
		#02 { a, b } = 8'b10100110;
		#02 { a, b } = 8'b10100111;
		#02 { a, b } = 8'b10101000;
		#02 { a, b } = 8'b10101001;
		#02 { a, b } = 8'b10101010;
		#02 { a, b } = 8'b10101011;
		#02 { a, b } = 8'b10101100;
		#02 { a, b } = 8'b10101101;
		#02 { a, b } = 8'b10101110;
		#02 { a, b } = 8'b10101111;
		#02 { a, b } = 8'b10110000;
		#02 { a, b } = 8'b10110001;
		#02 { a, b } = 8'b10110010;
		#02 { a, b } = 8'b10110011;
		#02 { a, b } = 8'b10110100;
		#02 { a, b } = 8'b10110101;
		#02 { a, b } = 8'b10110110;
		#02 { a, b } = 8'b10110111;
		#02 { a, b } = 8'b10111000;
		#02 { a, b } = 8'b10111001;
		#02 { a, b } = 8'b10111010;
		#02 { a, b } = 8'b10111011;
		#02 { a, b } = 8'b10111100;
		#02 { a, b } = 8'b10111101;
		#02 { a, b } = 8'b10111110;
		#02 { a, b } = 8'b10111111;
		#02 { a, b } = 8'b11000000;
		#02 { a, b } = 8'b11000001;
		#02 { a, b } = 8'b11000010;
		#02 { a, b } = 8'b11000011;
		#02 { a, b } = 8'b11000100;
		#02 { a, b } = 8'b11000101;
		#02 { a, b } = 8'b11000110;
		#02 { a, b } = 8'b11000111;
		#02 { a, b } = 8'b11001000;
		#02 { a, b } = 8'b11001001;
		#02 { a, b } = 8'b11001010;
		#02 { a, b } = 8'b11001011;
		#02 { a, b } = 8'b11001100;
		#02 { a, b } = 8'b11001101;
		#02 { a, b } = 8'b11001110;
		#02 { a, b } = 8'b11001111;
		#02 { a, b } = 8'b11010000;
		#02 { a, b } = 8'b11010001;
		#02 { a, b } = 8'b11010010;
		#02 { a, b } = 8'b11010011;
		#02 { a, b } = 8'b11010100;
		#02 { a, b } = 8'b11010101;
		#02 { a, b } = 8'b11010110;
		#02 { a, b } = 8'b11010111;
		#02 { a, b } = 8'b11011000;
		#02 { a, b } = 8'b11011001;
		#02 { a, b } = 8'b11011010;
		#02 { a, b } = 8'b11011011;
		#02 { a, b } = 8'b11011100;
		#02 { a, b } = 8'b11011101;
		#02 { a, b } = 8'b11011110;
		#02 { a, b } = 8'b11011111;
		#02 { a, b } = 8'b11100000;
		#02 { a, b } = 8'b11100001;
		#02 { a, b } = 8'b11100010;
		#02 { a, b } = 8'b11100011;
		#02 { a, b } = 8'b11100100;
		#02 { a, b } = 8'b11100101;
		#02 { a, b } = 8'b11100110;
		#02 { a, b } = 8'b11100111;
		#02 { a, b } = 8'b11101000;
		#02 { a, b } = 8'b11101001;
		#02 { a, b } = 8'b11101010;
		#02 { a, b } = 8'b11101011;
		#02 { a, b } = 8'b11101100;
		#02 { a, b } = 8'b11101101;
		#02 { a, b } = 8'b11101110;
		#02 { a, b } = 8'b11101111;
		#02 { a, b } = 8'b11110000;
		#02 { a, b } = 8'b11110001;
		#02 { a, b } = 8'b11110010;
		#02 { a, b } = 8'b11110011;
		#02 { a, b } = 8'b11110100;
		#02 { a, b } = 8'b11110101;
		#02 { a, b } = 8'b11110110;
		#02 { a, b } = 8'b11110111;
		#02 { a, b } = 8'b11111000;
		#02 { a, b } = 8'b11111001;
		#02 { a, b } = 8'b11111010;
		#02 { a, b } = 8'b11111011;
		#02 { a, b } = 8'b11111100;
		#02 { a, b } = 8'b11111101;
		#02 { a, b } = 8'b11111110;
		#02 { a, b } = 8'b11111111;
		#02 $finish;
	end
endmodule

module WorkBench;
	wire c;
	wire [3:0] a, b, s;
	TestGen test(s, c, a, b);
	Adder4b add(s, c, a, b);
endmodule
