/**
 * RISC: DMem.v
 * Author: Progyan Bhattacharya <progyanb@acm.org>
 *
 * This file contain Data Memory module. A Main Memory segment holding
 * 32-bit Data that has to be fetched by address.
 * A Test Generator module has been added for unit testing as well.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy of
 * this software and associated documentation files (the "Software"), to deal in
 * the Software without restriction, including without limitation the rights to use,
 * copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the
 * Software, and to permit persons to whom the Software is furnished to do so,
 * subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED,
 * INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A
 * PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF
 * CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE
 * OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 */

// Data Memory module
module DMem (
    output reg [31:0] rdata,
    input      [31:0] wdata, addr,
    input             clk, cnt);

    reg [31:0] dmem [0:1023];
    integer i;
    initial begin
        for ( i = 0; i < 1024; i = i + 1 )
            dmem[i] = 32'd0;
    end
    always @ ( negedge clk ) begin
        if ( cnt ) begin
            dmem[addr[9:0]] <= wdata;
            rdata <= wdata;
        end
        else
            rdata <= dmem[addr[9:0]];
    end
endmodule // DMem

// Test Generator Module to Test 1024x32-bit Data Memory
module TestDMem (
    input      [31:0] rdata,
    output reg [31:0] wdata, addr,
    input             clk,
    output reg        cnt);

    initial begin
        $monitor($time,,, "\nCC: %b\nAddress: %b\nData: %b\n", clk, addr, rdata);
            { cnt, addr } = { 1'b1, 10'd0 };
        #02 { cnt, addr } = { 1'b1, 10'd1 };
        #02 { cnt, addr } = { 1'b1, 10'd2 };
        #02 { cnt, addr } = { 1'b1, 10'd3 };
        #02 { cnt, addr } = { 1'b1, 10'd4 };
        #02 { cnt, addr } = { 1'b1, 10'd5 };
        #02 { cnt, addr } = { 1'b1, 10'd6 };
        #02 { cnt, addr } = { 1'b1, 10'd7 };
        #02 { cnt, addr } = { 1'b1, 10'd8 };
        #02 { cnt, addr } = { 1'b1, 10'd9 };
        #02 { cnt, addr } = { 1'b1, 10'd10 };
        #02 { cnt, addr } = { 1'b1, 10'd11 };
        #02 { cnt, addr } = { 1'b1, 10'd12 };
        #02 { cnt, addr } = { 1'b1, 10'd13 };
        #02 { cnt, addr } = { 1'b1, 10'd14 };
        #02 { cnt, addr } = { 1'b1, 10'd15 };
        #02 { cnt, addr } = { 1'b1, 10'd16 };
        #02 { cnt, addr } = { 1'b1, 10'd17 };
        #02 { cnt, addr } = { 1'b1, 10'd18 };
        #02 { cnt, addr } = { 1'b1, 10'd19 };
        #02 { cnt, addr } = { 1'b1, 10'd20 };
        #02 { cnt, addr } = { 1'b1, 10'd21 };
        #02 { cnt, addr } = { 1'b1, 10'd22 };
        #02 { cnt, addr } = { 1'b1, 10'd23 };
        #02 { cnt, addr } = { 1'b1, 10'd24 };
        #02 { cnt, addr } = { 1'b1, 10'd25 };
        #02 { cnt, addr } = { 1'b1, 10'd26 };
        #02 { cnt, addr } = { 1'b1, 10'd27 };
        #02 { cnt, addr } = { 1'b1, 10'd28 };
        #02 { cnt, addr } = { 1'b1, 10'd29 };
        #02 { cnt, addr } = { 1'b1, 10'd30 };
        #02 { cnt, addr } = { 1'b1, 10'd31 };
        #02 { cnt, addr } = { 1'b1, 10'd32 };
        #02 { cnt, addr } = { 1'b1, 10'd33 };
        #02 { cnt, addr } = { 1'b1, 10'd34 };
        #02 { cnt, addr } = { 1'b1, 10'd35 };
        #02 { cnt, addr } = { 1'b1, 10'd36 };
        #02 { cnt, addr } = { 1'b1, 10'd37 };
        #02 { cnt, addr } = { 1'b1, 10'd38 };
        #02 { cnt, addr } = { 1'b1, 10'd39 };
        #02 { cnt, addr } = { 1'b1, 10'd40 };
        #02 { cnt, addr } = { 1'b1, 10'd41 };
        #02 { cnt, addr } = { 1'b1, 10'd42 };
        #02 { cnt, addr } = { 1'b1, 10'd43 };
        #02 { cnt, addr } = { 1'b1, 10'd44 };
        #02 { cnt, addr } = { 1'b1, 10'd45 };
        #02 { cnt, addr } = { 1'b1, 10'd46 };
        #02 { cnt, addr } = { 1'b1, 10'd47 };
        #02 { cnt, addr } = { 1'b1, 10'd48 };
        #02 { cnt, addr } = { 1'b1, 10'd49 };
        #02 { cnt, addr } = { 1'b1, 10'd50 };
        #02 { cnt, addr } = { 1'b1, 10'd51 };
        #02 { cnt, addr } = { 1'b1, 10'd52 };
        #02 { cnt, addr } = { 1'b1, 10'd53 };
        #02 { cnt, addr } = { 1'b1, 10'd54 };
        #02 { cnt, addr } = { 1'b1, 10'd55 };
        #02 { cnt, addr } = { 1'b1, 10'd56 };
        #02 { cnt, addr } = { 1'b1, 10'd57 };
        #02 { cnt, addr } = { 1'b1, 10'd58 };
        #02 { cnt, addr } = { 1'b1, 10'd59 };
        #02 { cnt, addr } = { 1'b1, 10'd60 };
        #02 { cnt, addr } = { 1'b1, 10'd61 };
        #02 { cnt, addr } = { 1'b1, 10'd62 };
        #02 { cnt, addr } = { 1'b1, 10'd63 };
        #02 { cnt, addr } = { 1'b1, 10'd64 };
        #02 { cnt, addr } = { 1'b1, 10'd65 };
        #02 { cnt, addr } = { 1'b1, 10'd66 };
        #02 { cnt, addr } = { 1'b1, 10'd67 };
        #02 { cnt, addr } = { 1'b1, 10'd68 };
        #02 { cnt, addr } = { 1'b1, 10'd69 };
        #02 { cnt, addr } = { 1'b1, 10'd70 };
        #02 { cnt, addr } = { 1'b1, 10'd71 };
        #02 { cnt, addr } = { 1'b1, 10'd72 };
        #02 { cnt, addr } = { 1'b1, 10'd73 };
        #02 { cnt, addr } = { 1'b1, 10'd74 };
        #02 { cnt, addr } = { 1'b1, 10'd75 };
        #02 { cnt, addr } = { 1'b1, 10'd76 };
        #02 { cnt, addr } = { 1'b1, 10'd77 };
        #02 { cnt, addr } = { 1'b1, 10'd78 };
        #02 { cnt, addr } = { 1'b1, 10'd79 };
        #02 { cnt, addr } = { 1'b1, 10'd80 };
        #02 { cnt, addr } = { 1'b1, 10'd81 };
        #02 { cnt, addr } = { 1'b1, 10'd82 };
        #02 { cnt, addr } = { 1'b1, 10'd83 };
        #02 { cnt, addr } = { 1'b1, 10'd84 };
        #02 { cnt, addr } = { 1'b1, 10'd85 };
        #02 { cnt, addr } = { 1'b1, 10'd86 };
        #02 { cnt, addr } = { 1'b1, 10'd87 };
        #02 { cnt, addr } = { 1'b1, 10'd88 };
        #02 { cnt, addr } = { 1'b1, 10'd89 };
        #02 { cnt, addr } = { 1'b1, 10'd90 };
        #02 { cnt, addr } = { 1'b1, 10'd91 };
        #02 { cnt, addr } = { 1'b1, 10'd92 };
        #02 { cnt, addr } = { 1'b1, 10'd93 };
        #02 { cnt, addr } = { 1'b1, 10'd94 };
        #02 { cnt, addr } = { 1'b1, 10'd95 };
        #02 { cnt, addr } = { 1'b1, 10'd96 };
        #02 { cnt, addr } = { 1'b1, 10'd97 };
        #02 { cnt, addr } = { 1'b1, 10'd98 };
        #02 { cnt, addr } = { 1'b1, 10'd99 };
        #02 { cnt, addr } = { 1'b1, 10'd100 };
        #02 { cnt, addr } = { 1'b1, 10'd101 };
        #02 { cnt, addr } = { 1'b1, 10'd102 };
        #02 { cnt, addr } = { 1'b1, 10'd103 };
        #02 { cnt, addr } = { 1'b1, 10'd104 };
        #02 { cnt, addr } = { 1'b1, 10'd105 };
        #02 { cnt, addr } = { 1'b1, 10'd106 };
        #02 { cnt, addr } = { 1'b1, 10'd107 };
        #02 { cnt, addr } = { 1'b1, 10'd108 };
        #02 { cnt, addr } = { 1'b1, 10'd109 };
        #02 { cnt, addr } = { 1'b1, 10'd110 };
        #02 { cnt, addr } = { 1'b1, 10'd111 };
        #02 { cnt, addr } = { 1'b1, 10'd112 };
        #02 { cnt, addr } = { 1'b1, 10'd113 };
        #02 { cnt, addr } = { 1'b1, 10'd114 };
        #02 { cnt, addr } = { 1'b1, 10'd115 };
        #02 { cnt, addr } = { 1'b1, 10'd116 };
        #02 { cnt, addr } = { 1'b1, 10'd117 };
        #02 { cnt, addr } = { 1'b1, 10'd118 };
        #02 { cnt, addr } = { 1'b1, 10'd119 };
        #02 { cnt, addr } = { 1'b1, 10'd120 };
        #02 { cnt, addr } = { 1'b1, 10'd121 };
        #02 { cnt, addr } = { 1'b1, 10'd122 };
        #02 { cnt, addr } = { 1'b1, 10'd123 };
        #02 { cnt, addr } = { 1'b1, 10'd124 };
        #02 { cnt, addr } = { 1'b1, 10'd125 };
        #02 { cnt, addr } = { 1'b1, 10'd126 };
        #02 { cnt, addr } = { 1'b1, 10'd127 };
        #02 { cnt, addr } = { 1'b1, 10'd128 };
        #02 { cnt, addr } = { 1'b1, 10'd129 };
        #02 { cnt, addr } = { 1'b1, 10'd130 };
        #02 { cnt, addr } = { 1'b1, 10'd131 };
        #02 { cnt, addr } = { 1'b1, 10'd132 };
        #02 { cnt, addr } = { 1'b1, 10'd133 };
        #02 { cnt, addr } = { 1'b1, 10'd134 };
        #02 { cnt, addr } = { 1'b1, 10'd135 };
        #02 { cnt, addr } = { 1'b1, 10'd136 };
        #02 { cnt, addr } = { 1'b1, 10'd137 };
        #02 { cnt, addr } = { 1'b1, 10'd138 };
        #02 { cnt, addr } = { 1'b1, 10'd139 };
        #02 { cnt, addr } = { 1'b1, 10'd140 };
        #02 { cnt, addr } = { 1'b1, 10'd141 };
        #02 { cnt, addr } = { 1'b1, 10'd142 };
        #02 { cnt, addr } = { 1'b1, 10'd143 };
        #02 { cnt, addr } = { 1'b1, 10'd144 };
        #02 { cnt, addr } = { 1'b1, 10'd145 };
        #02 { cnt, addr } = { 1'b1, 10'd146 };
        #02 { cnt, addr } = { 1'b1, 10'd147 };
        #02 { cnt, addr } = { 1'b1, 10'd148 };
        #02 { cnt, addr } = { 1'b1, 10'd149 };
        #02 { cnt, addr } = { 1'b1, 10'd150 };
        #02 { cnt, addr } = { 1'b1, 10'd151 };
        #02 { cnt, addr } = { 1'b1, 10'd152 };
        #02 { cnt, addr } = { 1'b1, 10'd153 };
        #02 { cnt, addr } = { 1'b1, 10'd154 };
        #02 { cnt, addr } = { 1'b1, 10'd155 };
        #02 { cnt, addr } = { 1'b1, 10'd156 };
        #02 { cnt, addr } = { 1'b1, 10'd157 };
        #02 { cnt, addr } = { 1'b1, 10'd158 };
        #02 { cnt, addr } = { 1'b1, 10'd159 };
        #02 { cnt, addr } = { 1'b1, 10'd160 };
        #02 { cnt, addr } = { 1'b1, 10'd161 };
        #02 { cnt, addr } = { 1'b1, 10'd162 };
        #02 { cnt, addr } = { 1'b1, 10'd163 };
        #02 { cnt, addr } = { 1'b1, 10'd164 };
        #02 { cnt, addr } = { 1'b1, 10'd165 };
        #02 { cnt, addr } = { 1'b1, 10'd166 };
        #02 { cnt, addr } = { 1'b1, 10'd167 };
        #02 { cnt, addr } = { 1'b1, 10'd168 };
        #02 { cnt, addr } = { 1'b1, 10'd169 };
        #02 { cnt, addr } = { 1'b1, 10'd170 };
        #02 { cnt, addr } = { 1'b1, 10'd171 };
        #02 { cnt, addr } = { 1'b1, 10'd172 };
        #02 { cnt, addr } = { 1'b1, 10'd173 };
        #02 { cnt, addr } = { 1'b1, 10'd174 };
        #02 { cnt, addr } = { 1'b1, 10'd175 };
        #02 { cnt, addr } = { 1'b1, 10'd176 };
        #02 { cnt, addr } = { 1'b1, 10'd177 };
        #02 { cnt, addr } = { 1'b1, 10'd178 };
        #02 { cnt, addr } = { 1'b1, 10'd179 };
        #02 { cnt, addr } = { 1'b1, 10'd180 };
        #02 { cnt, addr } = { 1'b1, 10'd181 };
        #02 { cnt, addr } = { 1'b1, 10'd182 };
        #02 { cnt, addr } = { 1'b1, 10'd183 };
        #02 { cnt, addr } = { 1'b1, 10'd184 };
        #02 { cnt, addr } = { 1'b1, 10'd185 };
        #02 { cnt, addr } = { 1'b1, 10'd186 };
        #02 { cnt, addr } = { 1'b1, 10'd187 };
        #02 { cnt, addr } = { 1'b1, 10'd188 };
        #02 { cnt, addr } = { 1'b1, 10'd189 };
        #02 { cnt, addr } = { 1'b1, 10'd190 };
        #02 { cnt, addr } = { 1'b1, 10'd191 };
        #02 { cnt, addr } = { 1'b1, 10'd192 };
        #02 { cnt, addr } = { 1'b1, 10'd193 };
        #02 { cnt, addr } = { 1'b1, 10'd194 };
        #02 { cnt, addr } = { 1'b1, 10'd195 };
        #02 { cnt, addr } = { 1'b1, 10'd196 };
        #02 { cnt, addr } = { 1'b1, 10'd197 };
        #02 { cnt, addr } = { 1'b1, 10'd198 };
        #02 { cnt, addr } = { 1'b1, 10'd199 };
        #02 { cnt, addr } = { 1'b1, 10'd200 };
        #02 { cnt, addr } = { 1'b1, 10'd201 };
        #02 { cnt, addr } = { 1'b1, 10'd202 };
        #02 { cnt, addr } = { 1'b1, 10'd203 };
        #02 { cnt, addr } = { 1'b1, 10'd204 };
        #02 { cnt, addr } = { 1'b1, 10'd205 };
        #02 { cnt, addr } = { 1'b1, 10'd206 };
        #02 { cnt, addr } = { 1'b1, 10'd207 };
        #02 { cnt, addr } = { 1'b1, 10'd208 };
        #02 { cnt, addr } = { 1'b1, 10'd209 };
        #02 { cnt, addr } = { 1'b1, 10'd210 };
        #02 { cnt, addr } = { 1'b1, 10'd211 };
        #02 { cnt, addr } = { 1'b1, 10'd212 };
        #02 { cnt, addr } = { 1'b1, 10'd213 };
        #02 { cnt, addr } = { 1'b1, 10'd214 };
        #02 { cnt, addr } = { 1'b1, 10'd215 };
        #02 { cnt, addr } = { 1'b1, 10'd216 };
        #02 { cnt, addr } = { 1'b1, 10'd217 };
        #02 { cnt, addr } = { 1'b1, 10'd218 };
        #02 { cnt, addr } = { 1'b1, 10'd219 };
        #02 { cnt, addr } = { 1'b1, 10'd220 };
        #02 { cnt, addr } = { 1'b1, 10'd221 };
        #02 { cnt, addr } = { 1'b1, 10'd222 };
        #02 { cnt, addr } = { 1'b1, 10'd223 };
        #02 { cnt, addr } = { 1'b1, 10'd224 };
        #02 { cnt, addr } = { 1'b1, 10'd225 };
        #02 { cnt, addr } = { 1'b1, 10'd226 };
        #02 { cnt, addr } = { 1'b1, 10'd227 };
        #02 { cnt, addr } = { 1'b1, 10'd228 };
        #02 { cnt, addr } = { 1'b1, 10'd229 };
        #02 { cnt, addr } = { 1'b1, 10'd230 };
        #02 { cnt, addr } = { 1'b1, 10'd231 };
        #02 { cnt, addr } = { 1'b1, 10'd232 };
        #02 { cnt, addr } = { 1'b1, 10'd233 };
        #02 { cnt, addr } = { 1'b1, 10'd234 };
        #02 { cnt, addr } = { 1'b1, 10'd235 };
        #02 { cnt, addr } = { 1'b1, 10'd236 };
        #02 { cnt, addr } = { 1'b1, 10'd237 };
        #02 { cnt, addr } = { 1'b1, 10'd238 };
        #02 { cnt, addr } = { 1'b1, 10'd239 };
        #02 { cnt, addr } = { 1'b1, 10'd240 };
        #02 { cnt, addr } = { 1'b1, 10'd241 };
        #02 { cnt, addr } = { 1'b1, 10'd242 };
        #02 { cnt, addr } = { 1'b1, 10'd243 };
        #02 { cnt, addr } = { 1'b1, 10'd244 };
        #02 { cnt, addr } = { 1'b1, 10'd245 };
        #02 { cnt, addr } = { 1'b1, 10'd246 };
        #02 { cnt, addr } = { 1'b1, 10'd247 };
        #02 { cnt, addr } = { 1'b1, 10'd248 };
        #02 { cnt, addr } = { 1'b1, 10'd249 };
        #02 { cnt, addr } = { 1'b1, 10'd250 };
        #02 { cnt, addr } = { 1'b1, 10'd251 };
        #02 { cnt, addr } = { 1'b1, 10'd252 };
        #02 { cnt, addr } = { 1'b1, 10'd253 };
        #02 { cnt, addr } = { 1'b1, 10'd254 };
        #02 { cnt, addr } = { 1'b1, 10'd255 };
        #02 { cnt, addr } = { 1'b1, 10'd256 };
        #02 { cnt, addr } = { 1'b1, 10'd257 };
        #02 { cnt, addr } = { 1'b1, 10'd258 };
        #02 { cnt, addr } = { 1'b1, 10'd259 };
        #02 { cnt, addr } = { 1'b1, 10'd260 };
        #02 { cnt, addr } = { 1'b1, 10'd261 };
        #02 { cnt, addr } = { 1'b1, 10'd262 };
        #02 { cnt, addr } = { 1'b1, 10'd263 };
        #02 { cnt, addr } = { 1'b1, 10'd264 };
        #02 { cnt, addr } = { 1'b1, 10'd265 };
        #02 { cnt, addr } = { 1'b1, 10'd266 };
        #02 { cnt, addr } = { 1'b1, 10'd267 };
        #02 { cnt, addr } = { 1'b1, 10'd268 };
        #02 { cnt, addr } = { 1'b1, 10'd269 };
        #02 { cnt, addr } = { 1'b1, 10'd270 };
        #02 { cnt, addr } = { 1'b1, 10'd271 };
        #02 { cnt, addr } = { 1'b1, 10'd272 };
        #02 { cnt, addr } = { 1'b1, 10'd273 };
        #02 { cnt, addr } = { 1'b1, 10'd274 };
        #02 { cnt, addr } = { 1'b1, 10'd275 };
        #02 { cnt, addr } = { 1'b1, 10'd276 };
        #02 { cnt, addr } = { 1'b1, 10'd277 };
        #02 { cnt, addr } = { 1'b1, 10'd278 };
        #02 { cnt, addr } = { 1'b1, 10'd279 };
        #02 { cnt, addr } = { 1'b1, 10'd280 };
        #02 { cnt, addr } = { 1'b1, 10'd281 };
        #02 { cnt, addr } = { 1'b1, 10'd282 };
        #02 { cnt, addr } = { 1'b1, 10'd283 };
        #02 { cnt, addr } = { 1'b1, 10'd284 };
        #02 { cnt, addr } = { 1'b1, 10'd285 };
        #02 { cnt, addr } = { 1'b1, 10'd286 };
        #02 { cnt, addr } = { 1'b1, 10'd287 };
        #02 { cnt, addr } = { 1'b1, 10'd288 };
        #02 { cnt, addr } = { 1'b1, 10'd289 };
        #02 { cnt, addr } = { 1'b1, 10'd290 };
        #02 { cnt, addr } = { 1'b1, 10'd291 };
        #02 { cnt, addr } = { 1'b1, 10'd292 };
        #02 { cnt, addr } = { 1'b1, 10'd293 };
        #02 { cnt, addr } = { 1'b1, 10'd294 };
        #02 { cnt, addr } = { 1'b1, 10'd295 };
        #02 { cnt, addr } = { 1'b1, 10'd296 };
        #02 { cnt, addr } = { 1'b1, 10'd297 };
        #02 { cnt, addr } = { 1'b1, 10'd298 };
        #02 { cnt, addr } = { 1'b1, 10'd299 };
        #02 { cnt, addr } = { 1'b1, 10'd300 };
        #02 { cnt, addr } = { 1'b1, 10'd301 };
        #02 { cnt, addr } = { 1'b1, 10'd302 };
        #02 { cnt, addr } = { 1'b1, 10'd303 };
        #02 { cnt, addr } = { 1'b1, 10'd304 };
        #02 { cnt, addr } = { 1'b1, 10'd305 };
        #02 { cnt, addr } = { 1'b1, 10'd306 };
        #02 { cnt, addr } = { 1'b1, 10'd307 };
        #02 { cnt, addr } = { 1'b1, 10'd308 };
        #02 { cnt, addr } = { 1'b1, 10'd309 };
        #02 { cnt, addr } = { 1'b1, 10'd310 };
        #02 { cnt, addr } = { 1'b1, 10'd311 };
        #02 { cnt, addr } = { 1'b1, 10'd312 };
        #02 { cnt, addr } = { 1'b1, 10'd313 };
        #02 { cnt, addr } = { 1'b1, 10'd314 };
        #02 { cnt, addr } = { 1'b1, 10'd315 };
        #02 { cnt, addr } = { 1'b1, 10'd316 };
        #02 { cnt, addr } = { 1'b1, 10'd317 };
        #02 { cnt, addr } = { 1'b1, 10'd318 };
        #02 { cnt, addr } = { 1'b1, 10'd319 };
        #02 { cnt, addr } = { 1'b1, 10'd320 };
        #02 { cnt, addr } = { 1'b1, 10'd321 };
        #02 { cnt, addr } = { 1'b1, 10'd322 };
        #02 { cnt, addr } = { 1'b1, 10'd323 };
        #02 { cnt, addr } = { 1'b1, 10'd324 };
        #02 { cnt, addr } = { 1'b1, 10'd325 };
        #02 { cnt, addr } = { 1'b1, 10'd326 };
        #02 { cnt, addr } = { 1'b1, 10'd327 };
        #02 { cnt, addr } = { 1'b1, 10'd328 };
        #02 { cnt, addr } = { 1'b1, 10'd329 };
        #02 { cnt, addr } = { 1'b1, 10'd330 };
        #02 { cnt, addr } = { 1'b1, 10'd331 };
        #02 { cnt, addr } = { 1'b1, 10'd332 };
        #02 { cnt, addr } = { 1'b1, 10'd333 };
        #02 { cnt, addr } = { 1'b1, 10'd334 };
        #02 { cnt, addr } = { 1'b1, 10'd335 };
        #02 { cnt, addr } = { 1'b1, 10'd336 };
        #02 { cnt, addr } = { 1'b1, 10'd337 };
        #02 { cnt, addr } = { 1'b1, 10'd338 };
        #02 { cnt, addr } = { 1'b1, 10'd339 };
        #02 { cnt, addr } = { 1'b1, 10'd340 };
        #02 { cnt, addr } = { 1'b1, 10'd341 };
        #02 { cnt, addr } = { 1'b1, 10'd342 };
        #02 { cnt, addr } = { 1'b1, 10'd343 };
        #02 { cnt, addr } = { 1'b1, 10'd344 };
        #02 { cnt, addr } = { 1'b1, 10'd345 };
        #02 { cnt, addr } = { 1'b1, 10'd346 };
        #02 { cnt, addr } = { 1'b1, 10'd347 };
        #02 { cnt, addr } = { 1'b1, 10'd348 };
        #02 { cnt, addr } = { 1'b1, 10'd349 };
        #02 { cnt, addr } = { 1'b1, 10'd350 };
        #02 { cnt, addr } = { 1'b1, 10'd351 };
        #02 { cnt, addr } = { 1'b1, 10'd352 };
        #02 { cnt, addr } = { 1'b1, 10'd353 };
        #02 { cnt, addr } = { 1'b1, 10'd354 };
        #02 { cnt, addr } = { 1'b1, 10'd355 };
        #02 { cnt, addr } = { 1'b1, 10'd356 };
        #02 { cnt, addr } = { 1'b1, 10'd357 };
        #02 { cnt, addr } = { 1'b1, 10'd358 };
        #02 { cnt, addr } = { 1'b1, 10'd359 };
        #02 { cnt, addr } = { 1'b1, 10'd360 };
        #02 { cnt, addr } = { 1'b1, 10'd361 };
        #02 { cnt, addr } = { 1'b1, 10'd362 };
        #02 { cnt, addr } = { 1'b1, 10'd363 };
        #02 { cnt, addr } = { 1'b1, 10'd364 };
        #02 { cnt, addr } = { 1'b1, 10'd365 };
        #02 { cnt, addr } = { 1'b1, 10'd366 };
        #02 { cnt, addr } = { 1'b1, 10'd367 };
        #02 { cnt, addr } = { 1'b1, 10'd368 };
        #02 { cnt, addr } = { 1'b1, 10'd369 };
        #02 { cnt, addr } = { 1'b1, 10'd370 };
        #02 { cnt, addr } = { 1'b1, 10'd371 };
        #02 { cnt, addr } = { 1'b1, 10'd372 };
        #02 { cnt, addr } = { 1'b1, 10'd373 };
        #02 { cnt, addr } = { 1'b1, 10'd374 };
        #02 { cnt, addr } = { 1'b1, 10'd375 };
        #02 { cnt, addr } = { 1'b1, 10'd376 };
        #02 { cnt, addr } = { 1'b1, 10'd377 };
        #02 { cnt, addr } = { 1'b1, 10'd378 };
        #02 { cnt, addr } = { 1'b1, 10'd379 };
        #02 { cnt, addr } = { 1'b1, 10'd380 };
        #02 { cnt, addr } = { 1'b1, 10'd381 };
        #02 { cnt, addr } = { 1'b1, 10'd382 };
        #02 { cnt, addr } = { 1'b1, 10'd383 };
        #02 { cnt, addr } = { 1'b1, 10'd384 };
        #02 { cnt, addr } = { 1'b1, 10'd385 };
        #02 { cnt, addr } = { 1'b1, 10'd386 };
        #02 { cnt, addr } = { 1'b1, 10'd387 };
        #02 { cnt, addr } = { 1'b1, 10'd388 };
        #02 { cnt, addr } = { 1'b1, 10'd389 };
        #02 { cnt, addr } = { 1'b1, 10'd390 };
        #02 { cnt, addr } = { 1'b1, 10'd391 };
        #02 { cnt, addr } = { 1'b1, 10'd392 };
        #02 { cnt, addr } = { 1'b1, 10'd393 };
        #02 { cnt, addr } = { 1'b1, 10'd394 };
        #02 { cnt, addr } = { 1'b1, 10'd395 };
        #02 { cnt, addr } = { 1'b1, 10'd396 };
        #02 { cnt, addr } = { 1'b1, 10'd397 };
        #02 { cnt, addr } = { 1'b1, 10'd398 };
        #02 { cnt, addr } = { 1'b1, 10'd399 };
        #02 { cnt, addr } = { 1'b1, 10'd400 };
        #02 { cnt, addr } = { 1'b1, 10'd401 };
        #02 { cnt, addr } = { 1'b1, 10'd402 };
        #02 { cnt, addr } = { 1'b1, 10'd403 };
        #02 { cnt, addr } = { 1'b1, 10'd404 };
        #02 { cnt, addr } = { 1'b1, 10'd405 };
        #02 { cnt, addr } = { 1'b1, 10'd406 };
        #02 { cnt, addr } = { 1'b1, 10'd407 };
        #02 { cnt, addr } = { 1'b1, 10'd408 };
        #02 { cnt, addr } = { 1'b1, 10'd409 };
        #02 { cnt, addr } = { 1'b1, 10'd410 };
        #02 { cnt, addr } = { 1'b1, 10'd411 };
        #02 { cnt, addr } = { 1'b1, 10'd412 };
        #02 { cnt, addr } = { 1'b1, 10'd413 };
        #02 { cnt, addr } = { 1'b1, 10'd414 };
        #02 { cnt, addr } = { 1'b1, 10'd415 };
        #02 { cnt, addr } = { 1'b1, 10'd416 };
        #02 { cnt, addr } = { 1'b1, 10'd417 };
        #02 { cnt, addr } = { 1'b1, 10'd418 };
        #02 { cnt, addr } = { 1'b1, 10'd419 };
        #02 { cnt, addr } = { 1'b1, 10'd420 };
        #02 { cnt, addr } = { 1'b1, 10'd421 };
        #02 { cnt, addr } = { 1'b1, 10'd422 };
        #02 { cnt, addr } = { 1'b1, 10'd423 };
        #02 { cnt, addr } = { 1'b1, 10'd424 };
        #02 { cnt, addr } = { 1'b1, 10'd425 };
        #02 { cnt, addr } = { 1'b1, 10'd426 };
        #02 { cnt, addr } = { 1'b1, 10'd427 };
        #02 { cnt, addr } = { 1'b1, 10'd428 };
        #02 { cnt, addr } = { 1'b1, 10'd429 };
        #02 { cnt, addr } = { 1'b1, 10'd430 };
        #02 { cnt, addr } = { 1'b1, 10'd431 };
        #02 { cnt, addr } = { 1'b1, 10'd432 };
        #02 { cnt, addr } = { 1'b1, 10'd433 };
        #02 { cnt, addr } = { 1'b1, 10'd434 };
        #02 { cnt, addr } = { 1'b1, 10'd435 };
        #02 { cnt, addr } = { 1'b1, 10'd436 };
        #02 { cnt, addr } = { 1'b1, 10'd437 };
        #02 { cnt, addr } = { 1'b1, 10'd438 };
        #02 { cnt, addr } = { 1'b1, 10'd439 };
        #02 { cnt, addr } = { 1'b1, 10'd440 };
        #02 { cnt, addr } = { 1'b1, 10'd441 };
        #02 { cnt, addr } = { 1'b1, 10'd442 };
        #02 { cnt, addr } = { 1'b1, 10'd443 };
        #02 { cnt, addr } = { 1'b1, 10'd444 };
        #02 { cnt, addr } = { 1'b1, 10'd445 };
        #02 { cnt, addr } = { 1'b1, 10'd446 };
        #02 { cnt, addr } = { 1'b1, 10'd447 };
        #02 { cnt, addr } = { 1'b1, 10'd448 };
        #02 { cnt, addr } = { 1'b1, 10'd449 };
        #02 { cnt, addr } = { 1'b1, 10'd450 };
        #02 { cnt, addr } = { 1'b1, 10'd451 };
        #02 { cnt, addr } = { 1'b1, 10'd452 };
        #02 { cnt, addr } = { 1'b1, 10'd453 };
        #02 { cnt, addr } = { 1'b1, 10'd454 };
        #02 { cnt, addr } = { 1'b1, 10'd455 };
        #02 { cnt, addr } = { 1'b1, 10'd456 };
        #02 { cnt, addr } = { 1'b1, 10'd457 };
        #02 { cnt, addr } = { 1'b1, 10'd458 };
        #02 { cnt, addr } = { 1'b1, 10'd459 };
        #02 { cnt, addr } = { 1'b1, 10'd460 };
        #02 { cnt, addr } = { 1'b1, 10'd461 };
        #02 { cnt, addr } = { 1'b1, 10'd462 };
        #02 { cnt, addr } = { 1'b1, 10'd463 };
        #02 { cnt, addr } = { 1'b1, 10'd464 };
        #02 { cnt, addr } = { 1'b1, 10'd465 };
        #02 { cnt, addr } = { 1'b1, 10'd466 };
        #02 { cnt, addr } = { 1'b1, 10'd467 };
        #02 { cnt, addr } = { 1'b1, 10'd468 };
        #02 { cnt, addr } = { 1'b1, 10'd469 };
        #02 { cnt, addr } = { 1'b1, 10'd470 };
        #02 { cnt, addr } = { 1'b1, 10'd471 };
        #02 { cnt, addr } = { 1'b1, 10'd472 };
        #02 { cnt, addr } = { 1'b1, 10'd473 };
        #02 { cnt, addr } = { 1'b1, 10'd474 };
        #02 { cnt, addr } = { 1'b1, 10'd475 };
        #02 { cnt, addr } = { 1'b1, 10'd476 };
        #02 { cnt, addr } = { 1'b1, 10'd477 };
        #02 { cnt, addr } = { 1'b1, 10'd478 };
        #02 { cnt, addr } = { 1'b1, 10'd479 };
        #02 { cnt, addr } = { 1'b1, 10'd480 };
        #02 { cnt, addr } = { 1'b1, 10'd481 };
        #02 { cnt, addr } = { 1'b1, 10'd482 };
        #02 { cnt, addr } = { 1'b1, 10'd483 };
        #02 { cnt, addr } = { 1'b1, 10'd484 };
        #02 { cnt, addr } = { 1'b1, 10'd485 };
        #02 { cnt, addr } = { 1'b1, 10'd486 };
        #02 { cnt, addr } = { 1'b1, 10'd487 };
        #02 { cnt, addr } = { 1'b1, 10'd488 };
        #02 { cnt, addr } = { 1'b1, 10'd489 };
        #02 { cnt, addr } = { 1'b1, 10'd490 };
        #02 { cnt, addr } = { 1'b1, 10'd491 };
        #02 { cnt, addr } = { 1'b1, 10'd492 };
        #02 { cnt, addr } = { 1'b1, 10'd493 };
        #02 { cnt, addr } = { 1'b1, 10'd494 };
        #02 { cnt, addr } = { 1'b1, 10'd495 };
        #02 { cnt, addr } = { 1'b1, 10'd496 };
        #02 { cnt, addr } = { 1'b1, 10'd497 };
        #02 { cnt, addr } = { 1'b1, 10'd498 };
        #02 { cnt, addr } = { 1'b1, 10'd499 };
        #02 { cnt, addr } = { 1'b1, 10'd500 };
        #02 { cnt, addr } = { 1'b1, 10'd501 };
        #02 { cnt, addr } = { 1'b1, 10'd502 };
        #02 { cnt, addr } = { 1'b1, 10'd503 };
        #02 { cnt, addr } = { 1'b1, 10'd504 };
        #02 { cnt, addr } = { 1'b1, 10'd505 };
        #02 { cnt, addr } = { 1'b1, 10'd506 };
        #02 { cnt, addr } = { 1'b1, 10'd507 };
        #02 { cnt, addr } = { 1'b1, 10'd508 };
        #02 { cnt, addr } = { 1'b1, 10'd509 };
        #02 { cnt, addr } = { 1'b1, 10'd510 };
        #02 { cnt, addr } = { 1'b1, 10'd511 };
        #02 { cnt, addr } = { 1'b1, 10'd512 };
        #02 { cnt, addr } = { 1'b1, 10'd513 };
        #02 { cnt, addr } = { 1'b1, 10'd514 };
        #02 { cnt, addr } = { 1'b1, 10'd515 };
        #02 { cnt, addr } = { 1'b1, 10'd516 };
        #02 { cnt, addr } = { 1'b1, 10'd517 };
        #02 { cnt, addr } = { 1'b1, 10'd518 };
        #02 { cnt, addr } = { 1'b1, 10'd519 };
        #02 { cnt, addr } = { 1'b1, 10'd520 };
        #02 { cnt, addr } = { 1'b1, 10'd521 };
        #02 { cnt, addr } = { 1'b1, 10'd522 };
        #02 { cnt, addr } = { 1'b1, 10'd523 };
        #02 { cnt, addr } = { 1'b1, 10'd524 };
        #02 { cnt, addr } = { 1'b1, 10'd525 };
        #02 { cnt, addr } = { 1'b1, 10'd526 };
        #02 { cnt, addr } = { 1'b1, 10'd527 };
        #02 { cnt, addr } = { 1'b1, 10'd528 };
        #02 { cnt, addr } = { 1'b1, 10'd529 };
        #02 { cnt, addr } = { 1'b1, 10'd530 };
        #02 { cnt, addr } = { 1'b1, 10'd531 };
        #02 { cnt, addr } = { 1'b1, 10'd532 };
        #02 { cnt, addr } = { 1'b1, 10'd533 };
        #02 { cnt, addr } = { 1'b1, 10'd534 };
        #02 { cnt, addr } = { 1'b1, 10'd535 };
        #02 { cnt, addr } = { 1'b1, 10'd536 };
        #02 { cnt, addr } = { 1'b1, 10'd537 };
        #02 { cnt, addr } = { 1'b1, 10'd538 };
        #02 { cnt, addr } = { 1'b1, 10'd539 };
        #02 { cnt, addr } = { 1'b1, 10'd540 };
        #02 { cnt, addr } = { 1'b1, 10'd541 };
        #02 { cnt, addr } = { 1'b1, 10'd542 };
        #02 { cnt, addr } = { 1'b1, 10'd543 };
        #02 { cnt, addr } = { 1'b1, 10'd544 };
        #02 { cnt, addr } = { 1'b1, 10'd545 };
        #02 { cnt, addr } = { 1'b1, 10'd546 };
        #02 { cnt, addr } = { 1'b1, 10'd547 };
        #02 { cnt, addr } = { 1'b1, 10'd548 };
        #02 { cnt, addr } = { 1'b1, 10'd549 };
        #02 { cnt, addr } = { 1'b1, 10'd550 };
        #02 { cnt, addr } = { 1'b1, 10'd551 };
        #02 { cnt, addr } = { 1'b1, 10'd552 };
        #02 { cnt, addr } = { 1'b1, 10'd553 };
        #02 { cnt, addr } = { 1'b1, 10'd554 };
        #02 { cnt, addr } = { 1'b1, 10'd555 };
        #02 { cnt, addr } = { 1'b1, 10'd556 };
        #02 { cnt, addr } = { 1'b1, 10'd557 };
        #02 { cnt, addr } = { 1'b1, 10'd558 };
        #02 { cnt, addr } = { 1'b1, 10'd559 };
        #02 { cnt, addr } = { 1'b1, 10'd560 };
        #02 { cnt, addr } = { 1'b1, 10'd561 };
        #02 { cnt, addr } = { 1'b1, 10'd562 };
        #02 { cnt, addr } = { 1'b1, 10'd563 };
        #02 { cnt, addr } = { 1'b1, 10'd564 };
        #02 { cnt, addr } = { 1'b1, 10'd565 };
        #02 { cnt, addr } = { 1'b1, 10'd566 };
        #02 { cnt, addr } = { 1'b1, 10'd567 };
        #02 { cnt, addr } = { 1'b1, 10'd568 };
        #02 { cnt, addr } = { 1'b1, 10'd569 };
        #02 { cnt, addr } = { 1'b1, 10'd570 };
        #02 { cnt, addr } = { 1'b1, 10'd571 };
        #02 { cnt, addr } = { 1'b1, 10'd572 };
        #02 { cnt, addr } = { 1'b1, 10'd573 };
        #02 { cnt, addr } = { 1'b1, 10'd574 };
        #02 { cnt, addr } = { 1'b1, 10'd575 };
        #02 { cnt, addr } = { 1'b1, 10'd576 };
        #02 { cnt, addr } = { 1'b1, 10'd577 };
        #02 { cnt, addr } = { 1'b1, 10'd578 };
        #02 { cnt, addr } = { 1'b1, 10'd579 };
        #02 { cnt, addr } = { 1'b1, 10'd580 };
        #02 { cnt, addr } = { 1'b1, 10'd581 };
        #02 { cnt, addr } = { 1'b1, 10'd582 };
        #02 { cnt, addr } = { 1'b1, 10'd583 };
        #02 { cnt, addr } = { 1'b1, 10'd584 };
        #02 { cnt, addr } = { 1'b1, 10'd585 };
        #02 { cnt, addr } = { 1'b1, 10'd586 };
        #02 { cnt, addr } = { 1'b1, 10'd587 };
        #02 { cnt, addr } = { 1'b1, 10'd588 };
        #02 { cnt, addr } = { 1'b1, 10'd589 };
        #02 { cnt, addr } = { 1'b1, 10'd590 };
        #02 { cnt, addr } = { 1'b1, 10'd591 };
        #02 { cnt, addr } = { 1'b1, 10'd592 };
        #02 { cnt, addr } = { 1'b1, 10'd593 };
        #02 { cnt, addr } = { 1'b1, 10'd594 };
        #02 { cnt, addr } = { 1'b1, 10'd595 };
        #02 { cnt, addr } = { 1'b1, 10'd596 };
        #02 { cnt, addr } = { 1'b1, 10'd597 };
        #02 { cnt, addr } = { 1'b1, 10'd598 };
        #02 { cnt, addr } = { 1'b1, 10'd599 };
        #02 { cnt, addr } = { 1'b1, 10'd600 };
        #02 { cnt, addr } = { 1'b1, 10'd601 };
        #02 { cnt, addr } = { 1'b1, 10'd602 };
        #02 { cnt, addr } = { 1'b1, 10'd603 };
        #02 { cnt, addr } = { 1'b1, 10'd604 };
        #02 { cnt, addr } = { 1'b1, 10'd605 };
        #02 { cnt, addr } = { 1'b1, 10'd606 };
        #02 { cnt, addr } = { 1'b1, 10'd607 };
        #02 { cnt, addr } = { 1'b1, 10'd608 };
        #02 { cnt, addr } = { 1'b1, 10'd609 };
        #02 { cnt, addr } = { 1'b1, 10'd610 };
        #02 { cnt, addr } = { 1'b1, 10'd611 };
        #02 { cnt, addr } = { 1'b1, 10'd612 };
        #02 { cnt, addr } = { 1'b1, 10'd613 };
        #02 { cnt, addr } = { 1'b1, 10'd614 };
        #02 { cnt, addr } = { 1'b1, 10'd615 };
        #02 { cnt, addr } = { 1'b1, 10'd616 };
        #02 { cnt, addr } = { 1'b1, 10'd617 };
        #02 { cnt, addr } = { 1'b1, 10'd618 };
        #02 { cnt, addr } = { 1'b1, 10'd619 };
        #02 { cnt, addr } = { 1'b1, 10'd620 };
        #02 { cnt, addr } = { 1'b1, 10'd621 };
        #02 { cnt, addr } = { 1'b1, 10'd622 };
        #02 { cnt, addr } = { 1'b1, 10'd623 };
        #02 { cnt, addr } = { 1'b1, 10'd624 };
        #02 { cnt, addr } = { 1'b1, 10'd625 };
        #02 { cnt, addr } = { 1'b1, 10'd626 };
        #02 { cnt, addr } = { 1'b1, 10'd627 };
        #02 { cnt, addr } = { 1'b1, 10'd628 };
        #02 { cnt, addr } = { 1'b1, 10'd629 };
        #02 { cnt, addr } = { 1'b1, 10'd630 };
        #02 { cnt, addr } = { 1'b1, 10'd631 };
        #02 { cnt, addr } = { 1'b1, 10'd632 };
        #02 { cnt, addr } = { 1'b1, 10'd633 };
        #02 { cnt, addr } = { 1'b1, 10'd634 };
        #02 { cnt, addr } = { 1'b1, 10'd635 };
        #02 { cnt, addr } = { 1'b1, 10'd636 };
        #02 { cnt, addr } = { 1'b1, 10'd637 };
        #02 { cnt, addr } = { 1'b1, 10'd638 };
        #02 { cnt, addr } = { 1'b1, 10'd639 };
        #02 { cnt, addr } = { 1'b1, 10'd640 };
        #02 { cnt, addr } = { 1'b1, 10'd641 };
        #02 { cnt, addr } = { 1'b1, 10'd642 };
        #02 { cnt, addr } = { 1'b1, 10'd643 };
        #02 { cnt, addr } = { 1'b1, 10'd644 };
        #02 { cnt, addr } = { 1'b1, 10'd645 };
        #02 { cnt, addr } = { 1'b1, 10'd646 };
        #02 { cnt, addr } = { 1'b1, 10'd647 };
        #02 { cnt, addr } = { 1'b1, 10'd648 };
        #02 { cnt, addr } = { 1'b1, 10'd649 };
        #02 { cnt, addr } = { 1'b1, 10'd650 };
        #02 { cnt, addr } = { 1'b1, 10'd651 };
        #02 { cnt, addr } = { 1'b1, 10'd652 };
        #02 { cnt, addr } = { 1'b1, 10'd653 };
        #02 { cnt, addr } = { 1'b1, 10'd654 };
        #02 { cnt, addr } = { 1'b1, 10'd655 };
        #02 { cnt, addr } = { 1'b1, 10'd656 };
        #02 { cnt, addr } = { 1'b1, 10'd657 };
        #02 { cnt, addr } = { 1'b1, 10'd658 };
        #02 { cnt, addr } = { 1'b1, 10'd659 };
        #02 { cnt, addr } = { 1'b1, 10'd660 };
        #02 { cnt, addr } = { 1'b1, 10'd661 };
        #02 { cnt, addr } = { 1'b1, 10'd662 };
        #02 { cnt, addr } = { 1'b1, 10'd663 };
        #02 { cnt, addr } = { 1'b1, 10'd664 };
        #02 { cnt, addr } = { 1'b1, 10'd665 };
        #02 { cnt, addr } = { 1'b1, 10'd666 };
        #02 { cnt, addr } = { 1'b1, 10'd667 };
        #02 { cnt, addr } = { 1'b1, 10'd668 };
        #02 { cnt, addr } = { 1'b1, 10'd669 };
        #02 { cnt, addr } = { 1'b1, 10'd670 };
        #02 { cnt, addr } = { 1'b1, 10'd671 };
        #02 { cnt, addr } = { 1'b1, 10'd672 };
        #02 { cnt, addr } = { 1'b1, 10'd673 };
        #02 { cnt, addr } = { 1'b1, 10'd674 };
        #02 { cnt, addr } = { 1'b1, 10'd675 };
        #02 { cnt, addr } = { 1'b1, 10'd676 };
        #02 { cnt, addr } = { 1'b1, 10'd677 };
        #02 { cnt, addr } = { 1'b1, 10'd678 };
        #02 { cnt, addr } = { 1'b1, 10'd679 };
        #02 { cnt, addr } = { 1'b1, 10'd680 };
        #02 { cnt, addr } = { 1'b1, 10'd681 };
        #02 { cnt, addr } = { 1'b1, 10'd682 };
        #02 { cnt, addr } = { 1'b1, 10'd683 };
        #02 { cnt, addr } = { 1'b1, 10'd684 };
        #02 { cnt, addr } = { 1'b1, 10'd685 };
        #02 { cnt, addr } = { 1'b1, 10'd686 };
        #02 { cnt, addr } = { 1'b1, 10'd687 };
        #02 { cnt, addr } = { 1'b1, 10'd688 };
        #02 { cnt, addr } = { 1'b1, 10'd689 };
        #02 { cnt, addr } = { 1'b1, 10'd690 };
        #02 { cnt, addr } = { 1'b1, 10'd691 };
        #02 { cnt, addr } = { 1'b1, 10'd692 };
        #02 { cnt, addr } = { 1'b1, 10'd693 };
        #02 { cnt, addr } = { 1'b1, 10'd694 };
        #02 { cnt, addr } = { 1'b1, 10'd695 };
        #02 { cnt, addr } = { 1'b1, 10'd696 };
        #02 { cnt, addr } = { 1'b1, 10'd697 };
        #02 { cnt, addr } = { 1'b1, 10'd698 };
        #02 { cnt, addr } = { 1'b1, 10'd699 };
        #02 { cnt, addr } = { 1'b1, 10'd700 };
        #02 { cnt, addr } = { 1'b1, 10'd701 };
        #02 { cnt, addr } = { 1'b1, 10'd702 };
        #02 { cnt, addr } = { 1'b1, 10'd703 };
        #02 { cnt, addr } = { 1'b1, 10'd704 };
        #02 { cnt, addr } = { 1'b1, 10'd705 };
        #02 { cnt, addr } = { 1'b1, 10'd706 };
        #02 { cnt, addr } = { 1'b1, 10'd707 };
        #02 { cnt, addr } = { 1'b1, 10'd708 };
        #02 { cnt, addr } = { 1'b1, 10'd709 };
        #02 { cnt, addr } = { 1'b1, 10'd710 };
        #02 { cnt, addr } = { 1'b1, 10'd711 };
        #02 { cnt, addr } = { 1'b1, 10'd712 };
        #02 { cnt, addr } = { 1'b1, 10'd713 };
        #02 { cnt, addr } = { 1'b1, 10'd714 };
        #02 { cnt, addr } = { 1'b1, 10'd715 };
        #02 { cnt, addr } = { 1'b1, 10'd716 };
        #02 { cnt, addr } = { 1'b1, 10'd717 };
        #02 { cnt, addr } = { 1'b1, 10'd718 };
        #02 { cnt, addr } = { 1'b1, 10'd719 };
        #02 { cnt, addr } = { 1'b1, 10'd720 };
        #02 { cnt, addr } = { 1'b1, 10'd721 };
        #02 { cnt, addr } = { 1'b1, 10'd722 };
        #02 { cnt, addr } = { 1'b1, 10'd723 };
        #02 { cnt, addr } = { 1'b1, 10'd724 };
        #02 { cnt, addr } = { 1'b1, 10'd725 };
        #02 { cnt, addr } = { 1'b1, 10'd726 };
        #02 { cnt, addr } = { 1'b1, 10'd727 };
        #02 { cnt, addr } = { 1'b1, 10'd728 };
        #02 { cnt, addr } = { 1'b1, 10'd729 };
        #02 { cnt, addr } = { 1'b1, 10'd730 };
        #02 { cnt, addr } = { 1'b1, 10'd731 };
        #02 { cnt, addr } = { 1'b1, 10'd732 };
        #02 { cnt, addr } = { 1'b1, 10'd733 };
        #02 { cnt, addr } = { 1'b1, 10'd734 };
        #02 { cnt, addr } = { 1'b1, 10'd735 };
        #02 { cnt, addr } = { 1'b1, 10'd736 };
        #02 { cnt, addr } = { 1'b1, 10'd737 };
        #02 { cnt, addr } = { 1'b1, 10'd738 };
        #02 { cnt, addr } = { 1'b1, 10'd739 };
        #02 { cnt, addr } = { 1'b1, 10'd740 };
        #02 { cnt, addr } = { 1'b1, 10'd741 };
        #02 { cnt, addr } = { 1'b1, 10'd742 };
        #02 { cnt, addr } = { 1'b1, 10'd743 };
        #02 { cnt, addr } = { 1'b1, 10'd744 };
        #02 { cnt, addr } = { 1'b1, 10'd745 };
        #02 { cnt, addr } = { 1'b1, 10'd746 };
        #02 { cnt, addr } = { 1'b1, 10'd747 };
        #02 { cnt, addr } = { 1'b1, 10'd748 };
        #02 { cnt, addr } = { 1'b1, 10'd749 };
        #02 { cnt, addr } = { 1'b1, 10'd750 };
        #02 { cnt, addr } = { 1'b1, 10'd751 };
        #02 { cnt, addr } = { 1'b1, 10'd752 };
        #02 { cnt, addr } = { 1'b1, 10'd753 };
        #02 { cnt, addr } = { 1'b1, 10'd754 };
        #02 { cnt, addr } = { 1'b1, 10'd755 };
        #02 { cnt, addr } = { 1'b1, 10'd756 };
        #02 { cnt, addr } = { 1'b1, 10'd757 };
        #02 { cnt, addr } = { 1'b1, 10'd758 };
        #02 { cnt, addr } = { 1'b1, 10'd759 };
        #02 { cnt, addr } = { 1'b1, 10'd760 };
        #02 { cnt, addr } = { 1'b1, 10'd761 };
        #02 { cnt, addr } = { 1'b1, 10'd762 };
        #02 { cnt, addr } = { 1'b1, 10'd763 };
        #02 { cnt, addr } = { 1'b1, 10'd764 };
        #02 { cnt, addr } = { 1'b1, 10'd765 };
        #02 { cnt, addr } = { 1'b1, 10'd766 };
        #02 { cnt, addr } = { 1'b1, 10'd767 };
        #02 { cnt, addr } = { 1'b1, 10'd768 };
        #02 { cnt, addr } = { 1'b1, 10'd769 };
        #02 { cnt, addr } = { 1'b1, 10'd770 };
        #02 { cnt, addr } = { 1'b1, 10'd771 };
        #02 { cnt, addr } = { 1'b1, 10'd772 };
        #02 { cnt, addr } = { 1'b1, 10'd773 };
        #02 { cnt, addr } = { 1'b1, 10'd774 };
        #02 { cnt, addr } = { 1'b1, 10'd775 };
        #02 { cnt, addr } = { 1'b1, 10'd776 };
        #02 { cnt, addr } = { 1'b1, 10'd777 };
        #02 { cnt, addr } = { 1'b1, 10'd778 };
        #02 { cnt, addr } = { 1'b1, 10'd779 };
        #02 { cnt, addr } = { 1'b1, 10'd780 };
        #02 { cnt, addr } = { 1'b1, 10'd781 };
        #02 { cnt, addr } = { 1'b1, 10'd782 };
        #02 { cnt, addr } = { 1'b1, 10'd783 };
        #02 { cnt, addr } = { 1'b1, 10'd784 };
        #02 { cnt, addr } = { 1'b1, 10'd785 };
        #02 { cnt, addr } = { 1'b1, 10'd786 };
        #02 { cnt, addr } = { 1'b1, 10'd787 };
        #02 { cnt, addr } = { 1'b1, 10'd788 };
        #02 { cnt, addr } = { 1'b1, 10'd789 };
        #02 { cnt, addr } = { 1'b1, 10'd790 };
        #02 { cnt, addr } = { 1'b1, 10'd791 };
        #02 { cnt, addr } = { 1'b1, 10'd792 };
        #02 { cnt, addr } = { 1'b1, 10'd793 };
        #02 { cnt, addr } = { 1'b1, 10'd794 };
        #02 { cnt, addr } = { 1'b1, 10'd795 };
        #02 { cnt, addr } = { 1'b1, 10'd796 };
        #02 { cnt, addr } = { 1'b1, 10'd797 };
        #02 { cnt, addr } = { 1'b1, 10'd798 };
        #02 { cnt, addr } = { 1'b1, 10'd799 };
        #02 { cnt, addr } = { 1'b1, 10'd800 };
        #02 { cnt, addr } = { 1'b1, 10'd801 };
        #02 { cnt, addr } = { 1'b1, 10'd802 };
        #02 { cnt, addr } = { 1'b1, 10'd803 };
        #02 { cnt, addr } = { 1'b1, 10'd804 };
        #02 { cnt, addr } = { 1'b1, 10'd805 };
        #02 { cnt, addr } = { 1'b1, 10'd806 };
        #02 { cnt, addr } = { 1'b1, 10'd807 };
        #02 { cnt, addr } = { 1'b1, 10'd808 };
        #02 { cnt, addr } = { 1'b1, 10'd809 };
        #02 { cnt, addr } = { 1'b1, 10'd810 };
        #02 { cnt, addr } = { 1'b1, 10'd811 };
        #02 { cnt, addr } = { 1'b1, 10'd812 };
        #02 { cnt, addr } = { 1'b1, 10'd813 };
        #02 { cnt, addr } = { 1'b1, 10'd814 };
        #02 { cnt, addr } = { 1'b1, 10'd815 };
        #02 { cnt, addr } = { 1'b1, 10'd816 };
        #02 { cnt, addr } = { 1'b1, 10'd817 };
        #02 { cnt, addr } = { 1'b1, 10'd818 };
        #02 { cnt, addr } = { 1'b1, 10'd819 };
        #02 { cnt, addr } = { 1'b1, 10'd820 };
        #02 { cnt, addr } = { 1'b1, 10'd821 };
        #02 { cnt, addr } = { 1'b1, 10'd822 };
        #02 { cnt, addr } = { 1'b1, 10'd823 };
        #02 { cnt, addr } = { 1'b1, 10'd824 };
        #02 { cnt, addr } = { 1'b1, 10'd825 };
        #02 { cnt, addr } = { 1'b1, 10'd826 };
        #02 { cnt, addr } = { 1'b1, 10'd827 };
        #02 { cnt, addr } = { 1'b1, 10'd828 };
        #02 { cnt, addr } = { 1'b1, 10'd829 };
        #02 { cnt, addr } = { 1'b1, 10'd830 };
        #02 { cnt, addr } = { 1'b1, 10'd831 };
        #02 { cnt, addr } = { 1'b1, 10'd832 };
        #02 { cnt, addr } = { 1'b1, 10'd833 };
        #02 { cnt, addr } = { 1'b1, 10'd834 };
        #02 { cnt, addr } = { 1'b1, 10'd835 };
        #02 { cnt, addr } = { 1'b1, 10'd836 };
        #02 { cnt, addr } = { 1'b1, 10'd837 };
        #02 { cnt, addr } = { 1'b1, 10'd838 };
        #02 { cnt, addr } = { 1'b1, 10'd839 };
        #02 { cnt, addr } = { 1'b1, 10'd840 };
        #02 { cnt, addr } = { 1'b1, 10'd841 };
        #02 { cnt, addr } = { 1'b1, 10'd842 };
        #02 { cnt, addr } = { 1'b1, 10'd843 };
        #02 { cnt, addr } = { 1'b1, 10'd844 };
        #02 { cnt, addr } = { 1'b1, 10'd845 };
        #02 { cnt, addr } = { 1'b1, 10'd846 };
        #02 { cnt, addr } = { 1'b1, 10'd847 };
        #02 { cnt, addr } = { 1'b1, 10'd848 };
        #02 { cnt, addr } = { 1'b1, 10'd849 };
        #02 { cnt, addr } = { 1'b1, 10'd850 };
        #02 { cnt, addr } = { 1'b1, 10'd851 };
        #02 { cnt, addr } = { 1'b1, 10'd852 };
        #02 { cnt, addr } = { 1'b1, 10'd853 };
        #02 { cnt, addr } = { 1'b1, 10'd854 };
        #02 { cnt, addr } = { 1'b1, 10'd855 };
        #02 { cnt, addr } = { 1'b1, 10'd856 };
        #02 { cnt, addr } = { 1'b1, 10'd857 };
        #02 { cnt, addr } = { 1'b1, 10'd858 };
        #02 { cnt, addr } = { 1'b1, 10'd859 };
        #02 { cnt, addr } = { 1'b1, 10'd860 };
        #02 { cnt, addr } = { 1'b1, 10'd861 };
        #02 { cnt, addr } = { 1'b1, 10'd862 };
        #02 { cnt, addr } = { 1'b1, 10'd863 };
        #02 { cnt, addr } = { 1'b1, 10'd864 };
        #02 { cnt, addr } = { 1'b1, 10'd865 };
        #02 { cnt, addr } = { 1'b1, 10'd866 };
        #02 { cnt, addr } = { 1'b1, 10'd867 };
        #02 { cnt, addr } = { 1'b1, 10'd868 };
        #02 { cnt, addr } = { 1'b1, 10'd869 };
        #02 { cnt, addr } = { 1'b1, 10'd870 };
        #02 { cnt, addr } = { 1'b1, 10'd871 };
        #02 { cnt, addr } = { 1'b1, 10'd872 };
        #02 { cnt, addr } = { 1'b1, 10'd873 };
        #02 { cnt, addr } = { 1'b1, 10'd874 };
        #02 { cnt, addr } = { 1'b1, 10'd875 };
        #02 { cnt, addr } = { 1'b1, 10'd876 };
        #02 { cnt, addr } = { 1'b1, 10'd877 };
        #02 { cnt, addr } = { 1'b1, 10'd878 };
        #02 { cnt, addr } = { 1'b1, 10'd879 };
        #02 { cnt, addr } = { 1'b1, 10'd880 };
        #02 { cnt, addr } = { 1'b1, 10'd881 };
        #02 { cnt, addr } = { 1'b1, 10'd882 };
        #02 { cnt, addr } = { 1'b1, 10'd883 };
        #02 { cnt, addr } = { 1'b1, 10'd884 };
        #02 { cnt, addr } = { 1'b1, 10'd885 };
        #02 { cnt, addr } = { 1'b1, 10'd886 };
        #02 { cnt, addr } = { 1'b1, 10'd887 };
        #02 { cnt, addr } = { 1'b1, 10'd888 };
        #02 { cnt, addr } = { 1'b1, 10'd889 };
        #02 { cnt, addr } = { 1'b1, 10'd890 };
        #02 { cnt, addr } = { 1'b1, 10'd891 };
        #02 { cnt, addr } = { 1'b1, 10'd892 };
        #02 { cnt, addr } = { 1'b1, 10'd893 };
        #02 { cnt, addr } = { 1'b1, 10'd894 };
        #02 { cnt, addr } = { 1'b1, 10'd895 };
        #02 { cnt, addr } = { 1'b1, 10'd896 };
        #02 { cnt, addr } = { 1'b1, 10'd897 };
        #02 { cnt, addr } = { 1'b1, 10'd898 };
        #02 { cnt, addr } = { 1'b1, 10'd899 };
        #02 { cnt, addr } = { 1'b1, 10'd900 };
        #02 { cnt, addr } = { 1'b1, 10'd901 };
        #02 { cnt, addr } = { 1'b1, 10'd902 };
        #02 { cnt, addr } = { 1'b1, 10'd903 };
        #02 { cnt, addr } = { 1'b1, 10'd904 };
        #02 { cnt, addr } = { 1'b1, 10'd905 };
        #02 { cnt, addr } = { 1'b1, 10'd906 };
        #02 { cnt, addr } = { 1'b1, 10'd907 };
        #02 { cnt, addr } = { 1'b1, 10'd908 };
        #02 { cnt, addr } = { 1'b1, 10'd909 };
        #02 { cnt, addr } = { 1'b1, 10'd910 };
        #02 { cnt, addr } = { 1'b1, 10'd911 };
        #02 { cnt, addr } = { 1'b1, 10'd912 };
        #02 { cnt, addr } = { 1'b1, 10'd913 };
        #02 { cnt, addr } = { 1'b1, 10'd914 };
        #02 { cnt, addr } = { 1'b1, 10'd915 };
        #02 { cnt, addr } = { 1'b1, 10'd916 };
        #02 { cnt, addr } = { 1'b1, 10'd917 };
        #02 { cnt, addr } = { 1'b1, 10'd918 };
        #02 { cnt, addr } = { 1'b1, 10'd919 };
        #02 { cnt, addr } = { 1'b1, 10'd920 };
        #02 { cnt, addr } = { 1'b1, 10'd921 };
        #02 { cnt, addr } = { 1'b1, 10'd922 };
        #02 { cnt, addr } = { 1'b1, 10'd923 };
        #02 { cnt, addr } = { 1'b1, 10'd924 };
        #02 { cnt, addr } = { 1'b1, 10'd925 };
        #02 { cnt, addr } = { 1'b1, 10'd926 };
        #02 { cnt, addr } = { 1'b1, 10'd927 };
        #02 { cnt, addr } = { 1'b1, 10'd928 };
        #02 { cnt, addr } = { 1'b1, 10'd929 };
        #02 { cnt, addr } = { 1'b1, 10'd930 };
        #02 { cnt, addr } = { 1'b1, 10'd931 };
        #02 { cnt, addr } = { 1'b1, 10'd932 };
        #02 { cnt, addr } = { 1'b1, 10'd933 };
        #02 { cnt, addr } = { 1'b1, 10'd934 };
        #02 { cnt, addr } = { 1'b1, 10'd935 };
        #02 { cnt, addr } = { 1'b1, 10'd936 };
        #02 { cnt, addr } = { 1'b1, 10'd937 };
        #02 { cnt, addr } = { 1'b1, 10'd938 };
        #02 { cnt, addr } = { 1'b1, 10'd939 };
        #02 { cnt, addr } = { 1'b1, 10'd940 };
        #02 { cnt, addr } = { 1'b1, 10'd941 };
        #02 { cnt, addr } = { 1'b1, 10'd942 };
        #02 { cnt, addr } = { 1'b1, 10'd943 };
        #02 { cnt, addr } = { 1'b1, 10'd944 };
        #02 { cnt, addr } = { 1'b1, 10'd945 };
        #02 { cnt, addr } = { 1'b1, 10'd946 };
        #02 { cnt, addr } = { 1'b1, 10'd947 };
        #02 { cnt, addr } = { 1'b1, 10'd948 };
        #02 { cnt, addr } = { 1'b1, 10'd949 };
        #02 { cnt, addr } = { 1'b1, 10'd950 };
        #02 { cnt, addr } = { 1'b1, 10'd951 };
        #02 { cnt, addr } = { 1'b1, 10'd952 };
        #02 { cnt, addr } = { 1'b1, 10'd953 };
        #02 { cnt, addr } = { 1'b1, 10'd954 };
        #02 { cnt, addr } = { 1'b1, 10'd955 };
        #02 { cnt, addr } = { 1'b1, 10'd956 };
        #02 { cnt, addr } = { 1'b1, 10'd957 };
        #02 { cnt, addr } = { 1'b1, 10'd958 };
        #02 { cnt, addr } = { 1'b1, 10'd959 };
        #02 { cnt, addr } = { 1'b1, 10'd960 };
        #02 { cnt, addr } = { 1'b1, 10'd961 };
        #02 { cnt, addr } = { 1'b1, 10'd962 };
        #02 { cnt, addr } = { 1'b1, 10'd963 };
        #02 { cnt, addr } = { 1'b1, 10'd964 };
        #02 { cnt, addr } = { 1'b1, 10'd965 };
        #02 { cnt, addr } = { 1'b1, 10'd966 };
        #02 { cnt, addr } = { 1'b1, 10'd967 };
        #02 { cnt, addr } = { 1'b1, 10'd968 };
        #02 { cnt, addr } = { 1'b1, 10'd969 };
        #02 { cnt, addr } = { 1'b1, 10'd970 };
        #02 { cnt, addr } = { 1'b1, 10'd971 };
        #02 { cnt, addr } = { 1'b1, 10'd972 };
        #02 { cnt, addr } = { 1'b1, 10'd973 };
        #02 { cnt, addr } = { 1'b1, 10'd974 };
        #02 { cnt, addr } = { 1'b1, 10'd975 };
        #02 { cnt, addr } = { 1'b1, 10'd976 };
        #02 { cnt, addr } = { 1'b1, 10'd977 };
        #02 { cnt, addr } = { 1'b1, 10'd978 };
        #02 { cnt, addr } = { 1'b1, 10'd979 };
        #02 { cnt, addr } = { 1'b1, 10'd980 };
        #02 { cnt, addr } = { 1'b1, 10'd981 };
        #02 { cnt, addr } = { 1'b1, 10'd982 };
        #02 { cnt, addr } = { 1'b1, 10'd983 };
        #02 { cnt, addr } = { 1'b1, 10'd984 };
        #02 { cnt, addr } = { 1'b1, 10'd985 };
        #02 { cnt, addr } = { 1'b1, 10'd986 };
        #02 { cnt, addr } = { 1'b1, 10'd987 };
        #02 { cnt, addr } = { 1'b1, 10'd988 };
        #02 { cnt, addr } = { 1'b1, 10'd989 };
        #02 { cnt, addr } = { 1'b1, 10'd990 };
        #02 { cnt, addr } = { 1'b1, 10'd991 };
        #02 { cnt, addr } = { 1'b1, 10'd992 };
        #02 { cnt, addr } = { 1'b1, 10'd993 };
        #02 { cnt, addr } = { 1'b1, 10'd994 };
        #02 { cnt, addr } = { 1'b1, 10'd995 };
        #02 { cnt, addr } = { 1'b1, 10'd996 };
        #02 { cnt, addr } = { 1'b1, 10'd997 };
        #02 { cnt, addr } = { 1'b1, 10'd998 };
        #02 { cnt, addr } = { 1'b1, 10'd999 };
        #02 { cnt, addr } = { 1'b1, 10'd1000 };
        #02 { cnt, addr } = { 1'b1, 10'd1001 };
        #02 { cnt, addr } = { 1'b1, 10'd1002 };
        #02 { cnt, addr } = { 1'b1, 10'd1003 };
        #02 { cnt, addr } = { 1'b1, 10'd1004 };
        #02 { cnt, addr } = { 1'b1, 10'd1005 };
        #02 { cnt, addr } = { 1'b1, 10'd1006 };
        #02 { cnt, addr } = { 1'b1, 10'd1007 };
        #02 { cnt, addr } = { 1'b1, 10'd1008 };
        #02 { cnt, addr } = { 1'b1, 10'd1009 };
        #02 { cnt, addr } = { 1'b1, 10'd1010 };
        #02 { cnt, addr } = { 1'b1, 10'd1011 };
        #02 { cnt, addr } = { 1'b1, 10'd1012 };
        #02 { cnt, addr } = { 1'b1, 10'd1013 };
        #02 { cnt, addr } = { 1'b1, 10'd1014 };
        #02 { cnt, addr } = { 1'b1, 10'd1015 };
        #02 { cnt, addr } = { 1'b1, 10'd1016 };
        #02 { cnt, addr } = { 1'b1, 10'd1017 };
        #02 { cnt, addr } = { 1'b1, 10'd1018 };
        #02 { cnt, addr } = { 1'b1, 10'd1019 };
        #02 { cnt, addr } = { 1'b1, 10'd1020 };
        #02 { cnt, addr } = { 1'b1, 10'd1021 };
        #02 { cnt, addr } = { 1'b1, 10'd1022 };
        #02 { cnt, addr } = { 1'b1, 10'd1023 };
        #02 $finish;
    end
endmodule // TestDMem
