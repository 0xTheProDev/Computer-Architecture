/**
 * RISC: IMem.v
 * Author: Progyan Bhattacharya <progyanb@acm.org>
 *
 * This file contain Instruction Memory module. A Main Memory segment holding
 * 32-bit Instructions that has to be fetched by address.
 * A Test Generator module has been added for unit testing as well.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy of
 * this software and associated documentation files (the "Software"), to deal in
 * the Software without restriction, including without limitation the rights to use,
 * copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the
 * Software, and to permit persons to whom the Software is furnished to do so,
 * subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED,
 * INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A
 * PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
 * HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF
 * CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE
 * OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 */

// Instruction Memory module
module IMem (
    output reg [31:0] inst,
    input      [31:0] addr,
    input             clk);

    reg [31:0] imem [0:1023];
    // parameter ISource = "Instructions.txt";
    integer i;
    initial begin
        // $readmemh(ISource, imem, 0, 1023);
        for ( i = 0; i < 1024; i = i + 1 )
            imem[i] = 32'd0;
    end
    always @ ( * ) begin
        inst <= imem[addr[9:0]][31:0];
    end
endmodule // IMem

// Test Generator Module to Test 1024x32-bit Instruction Memory
module TestIMem (
    input      [31:0] inst,
    output reg [31:0] addr,
    input             clk);

    initial begin
        $monitor($time,,, "\nCC: %b\nAddress: %b\nInstruction: %b\n", clk, addr, inst);
            { addr } = { 10'd0 };
        #02 { addr } = { 10'd1 };
        #02 { addr } = { 10'd2 };
        #02 { addr } = { 10'd3 };
        #02 { addr } = { 10'd4 };
        #02 { addr } = { 10'd5 };
        #02 { addr } = { 10'd6 };
        #02 { addr } = { 10'd7 };
        #02 { addr } = { 10'd8 };
        #02 { addr } = { 10'd9 };
        #02 { addr } = { 10'd10 };
        #02 { addr } = { 10'd11 };
        #02 { addr } = { 10'd12 };
        #02 { addr } = { 10'd13 };
        #02 { addr } = { 10'd14 };
        #02 { addr } = { 10'd15 };
        #02 { addr } = { 10'd16 };
        #02 { addr } = { 10'd17 };
        #02 { addr } = { 10'd18 };
        #02 { addr } = { 10'd19 };
        #02 { addr } = { 10'd20 };
        #02 { addr } = { 10'd21 };
        #02 { addr } = { 10'd22 };
        #02 { addr } = { 10'd23 };
        #02 { addr } = { 10'd24 };
        #02 { addr } = { 10'd25 };
        #02 { addr } = { 10'd26 };
        #02 { addr } = { 10'd27 };
        #02 { addr } = { 10'd28 };
        #02 { addr } = { 10'd29 };
        #02 { addr } = { 10'd30 };
        #02 { addr } = { 10'd31 };
        #02 { addr } = { 10'd32 };
        #02 { addr } = { 10'd33 };
        #02 { addr } = { 10'd34 };
        #02 { addr } = { 10'd35 };
        #02 { addr } = { 10'd36 };
        #02 { addr } = { 10'd37 };
        #02 { addr } = { 10'd38 };
        #02 { addr } = { 10'd39 };
        #02 { addr } = { 10'd40 };
        #02 { addr } = { 10'd41 };
        #02 { addr } = { 10'd42 };
        #02 { addr } = { 10'd43 };
        #02 { addr } = { 10'd44 };
        #02 { addr } = { 10'd45 };
        #02 { addr } = { 10'd46 };
        #02 { addr } = { 10'd47 };
        #02 { addr } = { 10'd48 };
        #02 { addr } = { 10'd49 };
        #02 { addr } = { 10'd50 };
        #02 { addr } = { 10'd51 };
        #02 { addr } = { 10'd52 };
        #02 { addr } = { 10'd53 };
        #02 { addr } = { 10'd54 };
        #02 { addr } = { 10'd55 };
        #02 { addr } = { 10'd56 };
        #02 { addr } = { 10'd57 };
        #02 { addr } = { 10'd58 };
        #02 { addr } = { 10'd59 };
        #02 { addr } = { 10'd60 };
        #02 { addr } = { 10'd61 };
        #02 { addr } = { 10'd62 };
        #02 { addr } = { 10'd63 };
        #02 { addr } = { 10'd64 };
        #02 { addr } = { 10'd65 };
        #02 { addr } = { 10'd66 };
        #02 { addr } = { 10'd67 };
        #02 { addr } = { 10'd68 };
        #02 { addr } = { 10'd69 };
        #02 { addr } = { 10'd70 };
        #02 { addr } = { 10'd71 };
        #02 { addr } = { 10'd72 };
        #02 { addr } = { 10'd73 };
        #02 { addr } = { 10'd74 };
        #02 { addr } = { 10'd75 };
        #02 { addr } = { 10'd76 };
        #02 { addr } = { 10'd77 };
        #02 { addr } = { 10'd78 };
        #02 { addr } = { 10'd79 };
        #02 { addr } = { 10'd80 };
        #02 { addr } = { 10'd81 };
        #02 { addr } = { 10'd82 };
        #02 { addr } = { 10'd83 };
        #02 { addr } = { 10'd84 };
        #02 { addr } = { 10'd85 };
        #02 { addr } = { 10'd86 };
        #02 { addr } = { 10'd87 };
        #02 { addr } = { 10'd88 };
        #02 { addr } = { 10'd89 };
        #02 { addr } = { 10'd90 };
        #02 { addr } = { 10'd91 };
        #02 { addr } = { 10'd92 };
        #02 { addr } = { 10'd93 };
        #02 { addr } = { 10'd94 };
        #02 { addr } = { 10'd95 };
        #02 { addr } = { 10'd96 };
        #02 { addr } = { 10'd97 };
        #02 { addr } = { 10'd98 };
        #02 { addr } = { 10'd99 };
        #02 { addr } = { 10'd100 };
        #02 { addr } = { 10'd101 };
        #02 { addr } = { 10'd102 };
        #02 { addr } = { 10'd103 };
        #02 { addr } = { 10'd104 };
        #02 { addr } = { 10'd105 };
        #02 { addr } = { 10'd106 };
        #02 { addr } = { 10'd107 };
        #02 { addr } = { 10'd108 };
        #02 { addr } = { 10'd109 };
        #02 { addr } = { 10'd110 };
        #02 { addr } = { 10'd111 };
        #02 { addr } = { 10'd112 };
        #02 { addr } = { 10'd113 };
        #02 { addr } = { 10'd114 };
        #02 { addr } = { 10'd115 };
        #02 { addr } = { 10'd116 };
        #02 { addr } = { 10'd117 };
        #02 { addr } = { 10'd118 };
        #02 { addr } = { 10'd119 };
        #02 { addr } = { 10'd120 };
        #02 { addr } = { 10'd121 };
        #02 { addr } = { 10'd122 };
        #02 { addr } = { 10'd123 };
        #02 { addr } = { 10'd124 };
        #02 { addr } = { 10'd125 };
        #02 { addr } = { 10'd126 };
        #02 { addr } = { 10'd127 };
        #02 { addr } = { 10'd128 };
        #02 { addr } = { 10'd129 };
        #02 { addr } = { 10'd130 };
        #02 { addr } = { 10'd131 };
        #02 { addr } = { 10'd132 };
        #02 { addr } = { 10'd133 };
        #02 { addr } = { 10'd134 };
        #02 { addr } = { 10'd135 };
        #02 { addr } = { 10'd136 };
        #02 { addr } = { 10'd137 };
        #02 { addr } = { 10'd138 };
        #02 { addr } = { 10'd139 };
        #02 { addr } = { 10'd140 };
        #02 { addr } = { 10'd141 };
        #02 { addr } = { 10'd142 };
        #02 { addr } = { 10'd143 };
        #02 { addr } = { 10'd144 };
        #02 { addr } = { 10'd145 };
        #02 { addr } = { 10'd146 };
        #02 { addr } = { 10'd147 };
        #02 { addr } = { 10'd148 };
        #02 { addr } = { 10'd149 };
        #02 { addr } = { 10'd150 };
        #02 { addr } = { 10'd151 };
        #02 { addr } = { 10'd152 };
        #02 { addr } = { 10'd153 };
        #02 { addr } = { 10'd154 };
        #02 { addr } = { 10'd155 };
        #02 { addr } = { 10'd156 };
        #02 { addr } = { 10'd157 };
        #02 { addr } = { 10'd158 };
        #02 { addr } = { 10'd159 };
        #02 { addr } = { 10'd160 };
        #02 { addr } = { 10'd161 };
        #02 { addr } = { 10'd162 };
        #02 { addr } = { 10'd163 };
        #02 { addr } = { 10'd164 };
        #02 { addr } = { 10'd165 };
        #02 { addr } = { 10'd166 };
        #02 { addr } = { 10'd167 };
        #02 { addr } = { 10'd168 };
        #02 { addr } = { 10'd169 };
        #02 { addr } = { 10'd170 };
        #02 { addr } = { 10'd171 };
        #02 { addr } = { 10'd172 };
        #02 { addr } = { 10'd173 };
        #02 { addr } = { 10'd174 };
        #02 { addr } = { 10'd175 };
        #02 { addr } = { 10'd176 };
        #02 { addr } = { 10'd177 };
        #02 { addr } = { 10'd178 };
        #02 { addr } = { 10'd179 };
        #02 { addr } = { 10'd180 };
        #02 { addr } = { 10'd181 };
        #02 { addr } = { 10'd182 };
        #02 { addr } = { 10'd183 };
        #02 { addr } = { 10'd184 };
        #02 { addr } = { 10'd185 };
        #02 { addr } = { 10'd186 };
        #02 { addr } = { 10'd187 };
        #02 { addr } = { 10'd188 };
        #02 { addr } = { 10'd189 };
        #02 { addr } = { 10'd190 };
        #02 { addr } = { 10'd191 };
        #02 { addr } = { 10'd192 };
        #02 { addr } = { 10'd193 };
        #02 { addr } = { 10'd194 };
        #02 { addr } = { 10'd195 };
        #02 { addr } = { 10'd196 };
        #02 { addr } = { 10'd197 };
        #02 { addr } = { 10'd198 };
        #02 { addr } = { 10'd199 };
        #02 { addr } = { 10'd200 };
        #02 { addr } = { 10'd201 };
        #02 { addr } = { 10'd202 };
        #02 { addr } = { 10'd203 };
        #02 { addr } = { 10'd204 };
        #02 { addr } = { 10'd205 };
        #02 { addr } = { 10'd206 };
        #02 { addr } = { 10'd207 };
        #02 { addr } = { 10'd208 };
        #02 { addr } = { 10'd209 };
        #02 { addr } = { 10'd210 };
        #02 { addr } = { 10'd211 };
        #02 { addr } = { 10'd212 };
        #02 { addr } = { 10'd213 };
        #02 { addr } = { 10'd214 };
        #02 { addr } = { 10'd215 };
        #02 { addr } = { 10'd216 };
        #02 { addr } = { 10'd217 };
        #02 { addr } = { 10'd218 };
        #02 { addr } = { 10'd219 };
        #02 { addr } = { 10'd220 };
        #02 { addr } = { 10'd221 };
        #02 { addr } = { 10'd222 };
        #02 { addr } = { 10'd223 };
        #02 { addr } = { 10'd224 };
        #02 { addr } = { 10'd225 };
        #02 { addr } = { 10'd226 };
        #02 { addr } = { 10'd227 };
        #02 { addr } = { 10'd228 };
        #02 { addr } = { 10'd229 };
        #02 { addr } = { 10'd230 };
        #02 { addr } = { 10'd231 };
        #02 { addr } = { 10'd232 };
        #02 { addr } = { 10'd233 };
        #02 { addr } = { 10'd234 };
        #02 { addr } = { 10'd235 };
        #02 { addr } = { 10'd236 };
        #02 { addr } = { 10'd237 };
        #02 { addr } = { 10'd238 };
        #02 { addr } = { 10'd239 };
        #02 { addr } = { 10'd240 };
        #02 { addr } = { 10'd241 };
        #02 { addr } = { 10'd242 };
        #02 { addr } = { 10'd243 };
        #02 { addr } = { 10'd244 };
        #02 { addr } = { 10'd245 };
        #02 { addr } = { 10'd246 };
        #02 { addr } = { 10'd247 };
        #02 { addr } = { 10'd248 };
        #02 { addr } = { 10'd249 };
        #02 { addr } = { 10'd250 };
        #02 { addr } = { 10'd251 };
        #02 { addr } = { 10'd252 };
        #02 { addr } = { 10'd253 };
        #02 { addr } = { 10'd254 };
        #02 { addr } = { 10'd255 };
        #02 { addr } = { 10'd256 };
        #02 { addr } = { 10'd257 };
        #02 { addr } = { 10'd258 };
        #02 { addr } = { 10'd259 };
        #02 { addr } = { 10'd260 };
        #02 { addr } = { 10'd261 };
        #02 { addr } = { 10'd262 };
        #02 { addr } = { 10'd263 };
        #02 { addr } = { 10'd264 };
        #02 { addr } = { 10'd265 };
        #02 { addr } = { 10'd266 };
        #02 { addr } = { 10'd267 };
        #02 { addr } = { 10'd268 };
        #02 { addr } = { 10'd269 };
        #02 { addr } = { 10'd270 };
        #02 { addr } = { 10'd271 };
        #02 { addr } = { 10'd272 };
        #02 { addr } = { 10'd273 };
        #02 { addr } = { 10'd274 };
        #02 { addr } = { 10'd275 };
        #02 { addr } = { 10'd276 };
        #02 { addr } = { 10'd277 };
        #02 { addr } = { 10'd278 };
        #02 { addr } = { 10'd279 };
        #02 { addr } = { 10'd280 };
        #02 { addr } = { 10'd281 };
        #02 { addr } = { 10'd282 };
        #02 { addr } = { 10'd283 };
        #02 { addr } = { 10'd284 };
        #02 { addr } = { 10'd285 };
        #02 { addr } = { 10'd286 };
        #02 { addr } = { 10'd287 };
        #02 { addr } = { 10'd288 };
        #02 { addr } = { 10'd289 };
        #02 { addr } = { 10'd290 };
        #02 { addr } = { 10'd291 };
        #02 { addr } = { 10'd292 };
        #02 { addr } = { 10'd293 };
        #02 { addr } = { 10'd294 };
        #02 { addr } = { 10'd295 };
        #02 { addr } = { 10'd296 };
        #02 { addr } = { 10'd297 };
        #02 { addr } = { 10'd298 };
        #02 { addr } = { 10'd299 };
        #02 { addr } = { 10'd300 };
        #02 { addr } = { 10'd301 };
        #02 { addr } = { 10'd302 };
        #02 { addr } = { 10'd303 };
        #02 { addr } = { 10'd304 };
        #02 { addr } = { 10'd305 };
        #02 { addr } = { 10'd306 };
        #02 { addr } = { 10'd307 };
        #02 { addr } = { 10'd308 };
        #02 { addr } = { 10'd309 };
        #02 { addr } = { 10'd310 };
        #02 { addr } = { 10'd311 };
        #02 { addr } = { 10'd312 };
        #02 { addr } = { 10'd313 };
        #02 { addr } = { 10'd314 };
        #02 { addr } = { 10'd315 };
        #02 { addr } = { 10'd316 };
        #02 { addr } = { 10'd317 };
        #02 { addr } = { 10'd318 };
        #02 { addr } = { 10'd319 };
        #02 { addr } = { 10'd320 };
        #02 { addr } = { 10'd321 };
        #02 { addr } = { 10'd322 };
        #02 { addr } = { 10'd323 };
        #02 { addr } = { 10'd324 };
        #02 { addr } = { 10'd325 };
        #02 { addr } = { 10'd326 };
        #02 { addr } = { 10'd327 };
        #02 { addr } = { 10'd328 };
        #02 { addr } = { 10'd329 };
        #02 { addr } = { 10'd330 };
        #02 { addr } = { 10'd331 };
        #02 { addr } = { 10'd332 };
        #02 { addr } = { 10'd333 };
        #02 { addr } = { 10'd334 };
        #02 { addr } = { 10'd335 };
        #02 { addr } = { 10'd336 };
        #02 { addr } = { 10'd337 };
        #02 { addr } = { 10'd338 };
        #02 { addr } = { 10'd339 };
        #02 { addr } = { 10'd340 };
        #02 { addr } = { 10'd341 };
        #02 { addr } = { 10'd342 };
        #02 { addr } = { 10'd343 };
        #02 { addr } = { 10'd344 };
        #02 { addr } = { 10'd345 };
        #02 { addr } = { 10'd346 };
        #02 { addr } = { 10'd347 };
        #02 { addr } = { 10'd348 };
        #02 { addr } = { 10'd349 };
        #02 { addr } = { 10'd350 };
        #02 { addr } = { 10'd351 };
        #02 { addr } = { 10'd352 };
        #02 { addr } = { 10'd353 };
        #02 { addr } = { 10'd354 };
        #02 { addr } = { 10'd355 };
        #02 { addr } = { 10'd356 };
        #02 { addr } = { 10'd357 };
        #02 { addr } = { 10'd358 };
        #02 { addr } = { 10'd359 };
        #02 { addr } = { 10'd360 };
        #02 { addr } = { 10'd361 };
        #02 { addr } = { 10'd362 };
        #02 { addr } = { 10'd363 };
        #02 { addr } = { 10'd364 };
        #02 { addr } = { 10'd365 };
        #02 { addr } = { 10'd366 };
        #02 { addr } = { 10'd367 };
        #02 { addr } = { 10'd368 };
        #02 { addr } = { 10'd369 };
        #02 { addr } = { 10'd370 };
        #02 { addr } = { 10'd371 };
        #02 { addr } = { 10'd372 };
        #02 { addr } = { 10'd373 };
        #02 { addr } = { 10'd374 };
        #02 { addr } = { 10'd375 };
        #02 { addr } = { 10'd376 };
        #02 { addr } = { 10'd377 };
        #02 { addr } = { 10'd378 };
        #02 { addr } = { 10'd379 };
        #02 { addr } = { 10'd380 };
        #02 { addr } = { 10'd381 };
        #02 { addr } = { 10'd382 };
        #02 { addr } = { 10'd383 };
        #02 { addr } = { 10'd384 };
        #02 { addr } = { 10'd385 };
        #02 { addr } = { 10'd386 };
        #02 { addr } = { 10'd387 };
        #02 { addr } = { 10'd388 };
        #02 { addr } = { 10'd389 };
        #02 { addr } = { 10'd390 };
        #02 { addr } = { 10'd391 };
        #02 { addr } = { 10'd392 };
        #02 { addr } = { 10'd393 };
        #02 { addr } = { 10'd394 };
        #02 { addr } = { 10'd395 };
        #02 { addr } = { 10'd396 };
        #02 { addr } = { 10'd397 };
        #02 { addr } = { 10'd398 };
        #02 { addr } = { 10'd399 };
        #02 { addr } = { 10'd400 };
        #02 { addr } = { 10'd401 };
        #02 { addr } = { 10'd402 };
        #02 { addr } = { 10'd403 };
        #02 { addr } = { 10'd404 };
        #02 { addr } = { 10'd405 };
        #02 { addr } = { 10'd406 };
        #02 { addr } = { 10'd407 };
        #02 { addr } = { 10'd408 };
        #02 { addr } = { 10'd409 };
        #02 { addr } = { 10'd410 };
        #02 { addr } = { 10'd411 };
        #02 { addr } = { 10'd412 };
        #02 { addr } = { 10'd413 };
        #02 { addr } = { 10'd414 };
        #02 { addr } = { 10'd415 };
        #02 { addr } = { 10'd416 };
        #02 { addr } = { 10'd417 };
        #02 { addr } = { 10'd418 };
        #02 { addr } = { 10'd419 };
        #02 { addr } = { 10'd420 };
        #02 { addr } = { 10'd421 };
        #02 { addr } = { 10'd422 };
        #02 { addr } = { 10'd423 };
        #02 { addr } = { 10'd424 };
        #02 { addr } = { 10'd425 };
        #02 { addr } = { 10'd426 };
        #02 { addr } = { 10'd427 };
        #02 { addr } = { 10'd428 };
        #02 { addr } = { 10'd429 };
        #02 { addr } = { 10'd430 };
        #02 { addr } = { 10'd431 };
        #02 { addr } = { 10'd432 };
        #02 { addr } = { 10'd433 };
        #02 { addr } = { 10'd434 };
        #02 { addr } = { 10'd435 };
        #02 { addr } = { 10'd436 };
        #02 { addr } = { 10'd437 };
        #02 { addr } = { 10'd438 };
        #02 { addr } = { 10'd439 };
        #02 { addr } = { 10'd440 };
        #02 { addr } = { 10'd441 };
        #02 { addr } = { 10'd442 };
        #02 { addr } = { 10'd443 };
        #02 { addr } = { 10'd444 };
        #02 { addr } = { 10'd445 };
        #02 { addr } = { 10'd446 };
        #02 { addr } = { 10'd447 };
        #02 { addr } = { 10'd448 };
        #02 { addr } = { 10'd449 };
        #02 { addr } = { 10'd450 };
        #02 { addr } = { 10'd451 };
        #02 { addr } = { 10'd452 };
        #02 { addr } = { 10'd453 };
        #02 { addr } = { 10'd454 };
        #02 { addr } = { 10'd455 };
        #02 { addr } = { 10'd456 };
        #02 { addr } = { 10'd457 };
        #02 { addr } = { 10'd458 };
        #02 { addr } = { 10'd459 };
        #02 { addr } = { 10'd460 };
        #02 { addr } = { 10'd461 };
        #02 { addr } = { 10'd462 };
        #02 { addr } = { 10'd463 };
        #02 { addr } = { 10'd464 };
        #02 { addr } = { 10'd465 };
        #02 { addr } = { 10'd466 };
        #02 { addr } = { 10'd467 };
        #02 { addr } = { 10'd468 };
        #02 { addr } = { 10'd469 };
        #02 { addr } = { 10'd470 };
        #02 { addr } = { 10'd471 };
        #02 { addr } = { 10'd472 };
        #02 { addr } = { 10'd473 };
        #02 { addr } = { 10'd474 };
        #02 { addr } = { 10'd475 };
        #02 { addr } = { 10'd476 };
        #02 { addr } = { 10'd477 };
        #02 { addr } = { 10'd478 };
        #02 { addr } = { 10'd479 };
        #02 { addr } = { 10'd480 };
        #02 { addr } = { 10'd481 };
        #02 { addr } = { 10'd482 };
        #02 { addr } = { 10'd483 };
        #02 { addr } = { 10'd484 };
        #02 { addr } = { 10'd485 };
        #02 { addr } = { 10'd486 };
        #02 { addr } = { 10'd487 };
        #02 { addr } = { 10'd488 };
        #02 { addr } = { 10'd489 };
        #02 { addr } = { 10'd490 };
        #02 { addr } = { 10'd491 };
        #02 { addr } = { 10'd492 };
        #02 { addr } = { 10'd493 };
        #02 { addr } = { 10'd494 };
        #02 { addr } = { 10'd495 };
        #02 { addr } = { 10'd496 };
        #02 { addr } = { 10'd497 };
        #02 { addr } = { 10'd498 };
        #02 { addr } = { 10'd499 };
        #02 { addr } = { 10'd500 };
        #02 { addr } = { 10'd501 };
        #02 { addr } = { 10'd502 };
        #02 { addr } = { 10'd503 };
        #02 { addr } = { 10'd504 };
        #02 { addr } = { 10'd505 };
        #02 { addr } = { 10'd506 };
        #02 { addr } = { 10'd507 };
        #02 { addr } = { 10'd508 };
        #02 { addr } = { 10'd509 };
        #02 { addr } = { 10'd510 };
        #02 { addr } = { 10'd511 };
        #02 { addr } = { 10'd512 };
        #02 { addr } = { 10'd513 };
        #02 { addr } = { 10'd514 };
        #02 { addr } = { 10'd515 };
        #02 { addr } = { 10'd516 };
        #02 { addr } = { 10'd517 };
        #02 { addr } = { 10'd518 };
        #02 { addr } = { 10'd519 };
        #02 { addr } = { 10'd520 };
        #02 { addr } = { 10'd521 };
        #02 { addr } = { 10'd522 };
        #02 { addr } = { 10'd523 };
        #02 { addr } = { 10'd524 };
        #02 { addr } = { 10'd525 };
        #02 { addr } = { 10'd526 };
        #02 { addr } = { 10'd527 };
        #02 { addr } = { 10'd528 };
        #02 { addr } = { 10'd529 };
        #02 { addr } = { 10'd530 };
        #02 { addr } = { 10'd531 };
        #02 { addr } = { 10'd532 };
        #02 { addr } = { 10'd533 };
        #02 { addr } = { 10'd534 };
        #02 { addr } = { 10'd535 };
        #02 { addr } = { 10'd536 };
        #02 { addr } = { 10'd537 };
        #02 { addr } = { 10'd538 };
        #02 { addr } = { 10'd539 };
        #02 { addr } = { 10'd540 };
        #02 { addr } = { 10'd541 };
        #02 { addr } = { 10'd542 };
        #02 { addr } = { 10'd543 };
        #02 { addr } = { 10'd544 };
        #02 { addr } = { 10'd545 };
        #02 { addr } = { 10'd546 };
        #02 { addr } = { 10'd547 };
        #02 { addr } = { 10'd548 };
        #02 { addr } = { 10'd549 };
        #02 { addr } = { 10'd550 };
        #02 { addr } = { 10'd551 };
        #02 { addr } = { 10'd552 };
        #02 { addr } = { 10'd553 };
        #02 { addr } = { 10'd554 };
        #02 { addr } = { 10'd555 };
        #02 { addr } = { 10'd556 };
        #02 { addr } = { 10'd557 };
        #02 { addr } = { 10'd558 };
        #02 { addr } = { 10'd559 };
        #02 { addr } = { 10'd560 };
        #02 { addr } = { 10'd561 };
        #02 { addr } = { 10'd562 };
        #02 { addr } = { 10'd563 };
        #02 { addr } = { 10'd564 };
        #02 { addr } = { 10'd565 };
        #02 { addr } = { 10'd566 };
        #02 { addr } = { 10'd567 };
        #02 { addr } = { 10'd568 };
        #02 { addr } = { 10'd569 };
        #02 { addr } = { 10'd570 };
        #02 { addr } = { 10'd571 };
        #02 { addr } = { 10'd572 };
        #02 { addr } = { 10'd573 };
        #02 { addr } = { 10'd574 };
        #02 { addr } = { 10'd575 };
        #02 { addr } = { 10'd576 };
        #02 { addr } = { 10'd577 };
        #02 { addr } = { 10'd578 };
        #02 { addr } = { 10'd579 };
        #02 { addr } = { 10'd580 };
        #02 { addr } = { 10'd581 };
        #02 { addr } = { 10'd582 };
        #02 { addr } = { 10'd583 };
        #02 { addr } = { 10'd584 };
        #02 { addr } = { 10'd585 };
        #02 { addr } = { 10'd586 };
        #02 { addr } = { 10'd587 };
        #02 { addr } = { 10'd588 };
        #02 { addr } = { 10'd589 };
        #02 { addr } = { 10'd590 };
        #02 { addr } = { 10'd591 };
        #02 { addr } = { 10'd592 };
        #02 { addr } = { 10'd593 };
        #02 { addr } = { 10'd594 };
        #02 { addr } = { 10'd595 };
        #02 { addr } = { 10'd596 };
        #02 { addr } = { 10'd597 };
        #02 { addr } = { 10'd598 };
        #02 { addr } = { 10'd599 };
        #02 { addr } = { 10'd600 };
        #02 { addr } = { 10'd601 };
        #02 { addr } = { 10'd602 };
        #02 { addr } = { 10'd603 };
        #02 { addr } = { 10'd604 };
        #02 { addr } = { 10'd605 };
        #02 { addr } = { 10'd606 };
        #02 { addr } = { 10'd607 };
        #02 { addr } = { 10'd608 };
        #02 { addr } = { 10'd609 };
        #02 { addr } = { 10'd610 };
        #02 { addr } = { 10'd611 };
        #02 { addr } = { 10'd612 };
        #02 { addr } = { 10'd613 };
        #02 { addr } = { 10'd614 };
        #02 { addr } = { 10'd615 };
        #02 { addr } = { 10'd616 };
        #02 { addr } = { 10'd617 };
        #02 { addr } = { 10'd618 };
        #02 { addr } = { 10'd619 };
        #02 { addr } = { 10'd620 };
        #02 { addr } = { 10'd621 };
        #02 { addr } = { 10'd622 };
        #02 { addr } = { 10'd623 };
        #02 { addr } = { 10'd624 };
        #02 { addr } = { 10'd625 };
        #02 { addr } = { 10'd626 };
        #02 { addr } = { 10'd627 };
        #02 { addr } = { 10'd628 };
        #02 { addr } = { 10'd629 };
        #02 { addr } = { 10'd630 };
        #02 { addr } = { 10'd631 };
        #02 { addr } = { 10'd632 };
        #02 { addr } = { 10'd633 };
        #02 { addr } = { 10'd634 };
        #02 { addr } = { 10'd635 };
        #02 { addr } = { 10'd636 };
        #02 { addr } = { 10'd637 };
        #02 { addr } = { 10'd638 };
        #02 { addr } = { 10'd639 };
        #02 { addr } = { 10'd640 };
        #02 { addr } = { 10'd641 };
        #02 { addr } = { 10'd642 };
        #02 { addr } = { 10'd643 };
        #02 { addr } = { 10'd644 };
        #02 { addr } = { 10'd645 };
        #02 { addr } = { 10'd646 };
        #02 { addr } = { 10'd647 };
        #02 { addr } = { 10'd648 };
        #02 { addr } = { 10'd649 };
        #02 { addr } = { 10'd650 };
        #02 { addr } = { 10'd651 };
        #02 { addr } = { 10'd652 };
        #02 { addr } = { 10'd653 };
        #02 { addr } = { 10'd654 };
        #02 { addr } = { 10'd655 };
        #02 { addr } = { 10'd656 };
        #02 { addr } = { 10'd657 };
        #02 { addr } = { 10'd658 };
        #02 { addr } = { 10'd659 };
        #02 { addr } = { 10'd660 };
        #02 { addr } = { 10'd661 };
        #02 { addr } = { 10'd662 };
        #02 { addr } = { 10'd663 };
        #02 { addr } = { 10'd664 };
        #02 { addr } = { 10'd665 };
        #02 { addr } = { 10'd666 };
        #02 { addr } = { 10'd667 };
        #02 { addr } = { 10'd668 };
        #02 { addr } = { 10'd669 };
        #02 { addr } = { 10'd670 };
        #02 { addr } = { 10'd671 };
        #02 { addr } = { 10'd672 };
        #02 { addr } = { 10'd673 };
        #02 { addr } = { 10'd674 };
        #02 { addr } = { 10'd675 };
        #02 { addr } = { 10'd676 };
        #02 { addr } = { 10'd677 };
        #02 { addr } = { 10'd678 };
        #02 { addr } = { 10'd679 };
        #02 { addr } = { 10'd680 };
        #02 { addr } = { 10'd681 };
        #02 { addr } = { 10'd682 };
        #02 { addr } = { 10'd683 };
        #02 { addr } = { 10'd684 };
        #02 { addr } = { 10'd685 };
        #02 { addr } = { 10'd686 };
        #02 { addr } = { 10'd687 };
        #02 { addr } = { 10'd688 };
        #02 { addr } = { 10'd689 };
        #02 { addr } = { 10'd690 };
        #02 { addr } = { 10'd691 };
        #02 { addr } = { 10'd692 };
        #02 { addr } = { 10'd693 };
        #02 { addr } = { 10'd694 };
        #02 { addr } = { 10'd695 };
        #02 { addr } = { 10'd696 };
        #02 { addr } = { 10'd697 };
        #02 { addr } = { 10'd698 };
        #02 { addr } = { 10'd699 };
        #02 { addr } = { 10'd700 };
        #02 { addr } = { 10'd701 };
        #02 { addr } = { 10'd702 };
        #02 { addr } = { 10'd703 };
        #02 { addr } = { 10'd704 };
        #02 { addr } = { 10'd705 };
        #02 { addr } = { 10'd706 };
        #02 { addr } = { 10'd707 };
        #02 { addr } = { 10'd708 };
        #02 { addr } = { 10'd709 };
        #02 { addr } = { 10'd710 };
        #02 { addr } = { 10'd711 };
        #02 { addr } = { 10'd712 };
        #02 { addr } = { 10'd713 };
        #02 { addr } = { 10'd714 };
        #02 { addr } = { 10'd715 };
        #02 { addr } = { 10'd716 };
        #02 { addr } = { 10'd717 };
        #02 { addr } = { 10'd718 };
        #02 { addr } = { 10'd719 };
        #02 { addr } = { 10'd720 };
        #02 { addr } = { 10'd721 };
        #02 { addr } = { 10'd722 };
        #02 { addr } = { 10'd723 };
        #02 { addr } = { 10'd724 };
        #02 { addr } = { 10'd725 };
        #02 { addr } = { 10'd726 };
        #02 { addr } = { 10'd727 };
        #02 { addr } = { 10'd728 };
        #02 { addr } = { 10'd729 };
        #02 { addr } = { 10'd730 };
        #02 { addr } = { 10'd731 };
        #02 { addr } = { 10'd732 };
        #02 { addr } = { 10'd733 };
        #02 { addr } = { 10'd734 };
        #02 { addr } = { 10'd735 };
        #02 { addr } = { 10'd736 };
        #02 { addr } = { 10'd737 };
        #02 { addr } = { 10'd738 };
        #02 { addr } = { 10'd739 };
        #02 { addr } = { 10'd740 };
        #02 { addr } = { 10'd741 };
        #02 { addr } = { 10'd742 };
        #02 { addr } = { 10'd743 };
        #02 { addr } = { 10'd744 };
        #02 { addr } = { 10'd745 };
        #02 { addr } = { 10'd746 };
        #02 { addr } = { 10'd747 };
        #02 { addr } = { 10'd748 };
        #02 { addr } = { 10'd749 };
        #02 { addr } = { 10'd750 };
        #02 { addr } = { 10'd751 };
        #02 { addr } = { 10'd752 };
        #02 { addr } = { 10'd753 };
        #02 { addr } = { 10'd754 };
        #02 { addr } = { 10'd755 };
        #02 { addr } = { 10'd756 };
        #02 { addr } = { 10'd757 };
        #02 { addr } = { 10'd758 };
        #02 { addr } = { 10'd759 };
        #02 { addr } = { 10'd760 };
        #02 { addr } = { 10'd761 };
        #02 { addr } = { 10'd762 };
        #02 { addr } = { 10'd763 };
        #02 { addr } = { 10'd764 };
        #02 { addr } = { 10'd765 };
        #02 { addr } = { 10'd766 };
        #02 { addr } = { 10'd767 };
        #02 { addr } = { 10'd768 };
        #02 { addr } = { 10'd769 };
        #02 { addr } = { 10'd770 };
        #02 { addr } = { 10'd771 };
        #02 { addr } = { 10'd772 };
        #02 { addr } = { 10'd773 };
        #02 { addr } = { 10'd774 };
        #02 { addr } = { 10'd775 };
        #02 { addr } = { 10'd776 };
        #02 { addr } = { 10'd777 };
        #02 { addr } = { 10'd778 };
        #02 { addr } = { 10'd779 };
        #02 { addr } = { 10'd780 };
        #02 { addr } = { 10'd781 };
        #02 { addr } = { 10'd782 };
        #02 { addr } = { 10'd783 };
        #02 { addr } = { 10'd784 };
        #02 { addr } = { 10'd785 };
        #02 { addr } = { 10'd786 };
        #02 { addr } = { 10'd787 };
        #02 { addr } = { 10'd788 };
        #02 { addr } = { 10'd789 };
        #02 { addr } = { 10'd790 };
        #02 { addr } = { 10'd791 };
        #02 { addr } = { 10'd792 };
        #02 { addr } = { 10'd793 };
        #02 { addr } = { 10'd794 };
        #02 { addr } = { 10'd795 };
        #02 { addr } = { 10'd796 };
        #02 { addr } = { 10'd797 };
        #02 { addr } = { 10'd798 };
        #02 { addr } = { 10'd799 };
        #02 { addr } = { 10'd800 };
        #02 { addr } = { 10'd801 };
        #02 { addr } = { 10'd802 };
        #02 { addr } = { 10'd803 };
        #02 { addr } = { 10'd804 };
        #02 { addr } = { 10'd805 };
        #02 { addr } = { 10'd806 };
        #02 { addr } = { 10'd807 };
        #02 { addr } = { 10'd808 };
        #02 { addr } = { 10'd809 };
        #02 { addr } = { 10'd810 };
        #02 { addr } = { 10'd811 };
        #02 { addr } = { 10'd812 };
        #02 { addr } = { 10'd813 };
        #02 { addr } = { 10'd814 };
        #02 { addr } = { 10'd815 };
        #02 { addr } = { 10'd816 };
        #02 { addr } = { 10'd817 };
        #02 { addr } = { 10'd818 };
        #02 { addr } = { 10'd819 };
        #02 { addr } = { 10'd820 };
        #02 { addr } = { 10'd821 };
        #02 { addr } = { 10'd822 };
        #02 { addr } = { 10'd823 };
        #02 { addr } = { 10'd824 };
        #02 { addr } = { 10'd825 };
        #02 { addr } = { 10'd826 };
        #02 { addr } = { 10'd827 };
        #02 { addr } = { 10'd828 };
        #02 { addr } = { 10'd829 };
        #02 { addr } = { 10'd830 };
        #02 { addr } = { 10'd831 };
        #02 { addr } = { 10'd832 };
        #02 { addr } = { 10'd833 };
        #02 { addr } = { 10'd834 };
        #02 { addr } = { 10'd835 };
        #02 { addr } = { 10'd836 };
        #02 { addr } = { 10'd837 };
        #02 { addr } = { 10'd838 };
        #02 { addr } = { 10'd839 };
        #02 { addr } = { 10'd840 };
        #02 { addr } = { 10'd841 };
        #02 { addr } = { 10'd842 };
        #02 { addr } = { 10'd843 };
        #02 { addr } = { 10'd844 };
        #02 { addr } = { 10'd845 };
        #02 { addr } = { 10'd846 };
        #02 { addr } = { 10'd847 };
        #02 { addr } = { 10'd848 };
        #02 { addr } = { 10'd849 };
        #02 { addr } = { 10'd850 };
        #02 { addr } = { 10'd851 };
        #02 { addr } = { 10'd852 };
        #02 { addr } = { 10'd853 };
        #02 { addr } = { 10'd854 };
        #02 { addr } = { 10'd855 };
        #02 { addr } = { 10'd856 };
        #02 { addr } = { 10'd857 };
        #02 { addr } = { 10'd858 };
        #02 { addr } = { 10'd859 };
        #02 { addr } = { 10'd860 };
        #02 { addr } = { 10'd861 };
        #02 { addr } = { 10'd862 };
        #02 { addr } = { 10'd863 };
        #02 { addr } = { 10'd864 };
        #02 { addr } = { 10'd865 };
        #02 { addr } = { 10'd866 };
        #02 { addr } = { 10'd867 };
        #02 { addr } = { 10'd868 };
        #02 { addr } = { 10'd869 };
        #02 { addr } = { 10'd870 };
        #02 { addr } = { 10'd871 };
        #02 { addr } = { 10'd872 };
        #02 { addr } = { 10'd873 };
        #02 { addr } = { 10'd874 };
        #02 { addr } = { 10'd875 };
        #02 { addr } = { 10'd876 };
        #02 { addr } = { 10'd877 };
        #02 { addr } = { 10'd878 };
        #02 { addr } = { 10'd879 };
        #02 { addr } = { 10'd880 };
        #02 { addr } = { 10'd881 };
        #02 { addr } = { 10'd882 };
        #02 { addr } = { 10'd883 };
        #02 { addr } = { 10'd884 };
        #02 { addr } = { 10'd885 };
        #02 { addr } = { 10'd886 };
        #02 { addr } = { 10'd887 };
        #02 { addr } = { 10'd888 };
        #02 { addr } = { 10'd889 };
        #02 { addr } = { 10'd890 };
        #02 { addr } = { 10'd891 };
        #02 { addr } = { 10'd892 };
        #02 { addr } = { 10'd893 };
        #02 { addr } = { 10'd894 };
        #02 { addr } = { 10'd895 };
        #02 { addr } = { 10'd896 };
        #02 { addr } = { 10'd897 };
        #02 { addr } = { 10'd898 };
        #02 { addr } = { 10'd899 };
        #02 { addr } = { 10'd900 };
        #02 { addr } = { 10'd901 };
        #02 { addr } = { 10'd902 };
        #02 { addr } = { 10'd903 };
        #02 { addr } = { 10'd904 };
        #02 { addr } = { 10'd905 };
        #02 { addr } = { 10'd906 };
        #02 { addr } = { 10'd907 };
        #02 { addr } = { 10'd908 };
        #02 { addr } = { 10'd909 };
        #02 { addr } = { 10'd910 };
        #02 { addr } = { 10'd911 };
        #02 { addr } = { 10'd912 };
        #02 { addr } = { 10'd913 };
        #02 { addr } = { 10'd914 };
        #02 { addr } = { 10'd915 };
        #02 { addr } = { 10'd916 };
        #02 { addr } = { 10'd917 };
        #02 { addr } = { 10'd918 };
        #02 { addr } = { 10'd919 };
        #02 { addr } = { 10'd920 };
        #02 { addr } = { 10'd921 };
        #02 { addr } = { 10'd922 };
        #02 { addr } = { 10'd923 };
        #02 { addr } = { 10'd924 };
        #02 { addr } = { 10'd925 };
        #02 { addr } = { 10'd926 };
        #02 { addr } = { 10'd927 };
        #02 { addr } = { 10'd928 };
        #02 { addr } = { 10'd929 };
        #02 { addr } = { 10'd930 };
        #02 { addr } = { 10'd931 };
        #02 { addr } = { 10'd932 };
        #02 { addr } = { 10'd933 };
        #02 { addr } = { 10'd934 };
        #02 { addr } = { 10'd935 };
        #02 { addr } = { 10'd936 };
        #02 { addr } = { 10'd937 };
        #02 { addr } = { 10'd938 };
        #02 { addr } = { 10'd939 };
        #02 { addr } = { 10'd940 };
        #02 { addr } = { 10'd941 };
        #02 { addr } = { 10'd942 };
        #02 { addr } = { 10'd943 };
        #02 { addr } = { 10'd944 };
        #02 { addr } = { 10'd945 };
        #02 { addr } = { 10'd946 };
        #02 { addr } = { 10'd947 };
        #02 { addr } = { 10'd948 };
        #02 { addr } = { 10'd949 };
        #02 { addr } = { 10'd950 };
        #02 { addr } = { 10'd951 };
        #02 { addr } = { 10'd952 };
        #02 { addr } = { 10'd953 };
        #02 { addr } = { 10'd954 };
        #02 { addr } = { 10'd955 };
        #02 { addr } = { 10'd956 };
        #02 { addr } = { 10'd957 };
        #02 { addr } = { 10'd958 };
        #02 { addr } = { 10'd959 };
        #02 { addr } = { 10'd960 };
        #02 { addr } = { 10'd961 };
        #02 { addr } = { 10'd962 };
        #02 { addr } = { 10'd963 };
        #02 { addr } = { 10'd964 };
        #02 { addr } = { 10'd965 };
        #02 { addr } = { 10'd966 };
        #02 { addr } = { 10'd967 };
        #02 { addr } = { 10'd968 };
        #02 { addr } = { 10'd969 };
        #02 { addr } = { 10'd970 };
        #02 { addr } = { 10'd971 };
        #02 { addr } = { 10'd972 };
        #02 { addr } = { 10'd973 };
        #02 { addr } = { 10'd974 };
        #02 { addr } = { 10'd975 };
        #02 { addr } = { 10'd976 };
        #02 { addr } = { 10'd977 };
        #02 { addr } = { 10'd978 };
        #02 { addr } = { 10'd979 };
        #02 { addr } = { 10'd980 };
        #02 { addr } = { 10'd981 };
        #02 { addr } = { 10'd982 };
        #02 { addr } = { 10'd983 };
        #02 { addr } = { 10'd984 };
        #02 { addr } = { 10'd985 };
        #02 { addr } = { 10'd986 };
        #02 { addr } = { 10'd987 };
        #02 { addr } = { 10'd988 };
        #02 { addr } = { 10'd989 };
        #02 { addr } = { 10'd990 };
        #02 { addr } = { 10'd991 };
        #02 { addr } = { 10'd992 };
        #02 { addr } = { 10'd993 };
        #02 { addr } = { 10'd994 };
        #02 { addr } = { 10'd995 };
        #02 { addr } = { 10'd996 };
        #02 { addr } = { 10'd997 };
        #02 { addr } = { 10'd998 };
        #02 { addr } = { 10'd999 };
        #02 { addr } = { 10'd1000 };
        #02 { addr } = { 10'd1001 };
        #02 { addr } = { 10'd1002 };
        #02 { addr } = { 10'd1003 };
        #02 { addr } = { 10'd1004 };
        #02 { addr } = { 10'd1005 };
        #02 { addr } = { 10'd1006 };
        #02 { addr } = { 10'd1007 };
        #02 { addr } = { 10'd1008 };
        #02 { addr } = { 10'd1009 };
        #02 { addr } = { 10'd1010 };
        #02 { addr } = { 10'd1011 };
        #02 { addr } = { 10'd1012 };
        #02 { addr } = { 10'd1013 };
        #02 { addr } = { 10'd1014 };
        #02 { addr } = { 10'd1015 };
        #02 { addr } = { 10'd1016 };
        #02 { addr } = { 10'd1017 };
        #02 { addr } = { 10'd1018 };
        #02 { addr } = { 10'd1019 };
        #02 { addr } = { 10'd1020 };
        #02 { addr } = { 10'd1021 };
        #02 { addr } = { 10'd1022 };
        #02 { addr } = { 10'd1023 };
        #02 $finish;
    end
endmodule // TestIMem
